magic
tech sky130A
timestamp 1717243586
<< pwell >>
rect -139 -454 139 454
<< mvnmos >>
rect -25 -325 25 325
<< mvndiff >>
rect -54 319 -25 325
rect -54 -319 -48 319
rect -31 -319 -25 319
rect -54 -325 -25 -319
rect 25 319 54 325
rect 25 -319 31 319
rect 48 -319 54 319
rect 25 -325 54 -319
<< mvndiffc >>
rect -48 -319 -31 319
rect 31 -319 48 319
<< mvpsubdiff >>
rect -121 430 121 436
rect -121 413 -67 430
rect 67 413 121 430
rect -121 407 121 413
rect -121 382 -92 407
rect -121 -382 -115 382
rect -98 -382 -92 382
rect 92 382 121 407
rect -121 -407 -92 -382
rect 92 -382 98 382
rect 115 -382 121 382
rect 92 -407 121 -382
rect -121 -413 121 -407
rect -121 -430 -67 -413
rect 67 -430 121 -413
rect -121 -436 121 -430
<< mvpsubdiffcont >>
rect -67 413 67 430
rect -115 -382 -98 382
rect 98 -382 115 382
rect -67 -430 67 -413
<< poly >>
rect -25 361 25 369
rect -25 344 -17 361
rect 17 344 25 361
rect -25 325 25 344
rect -25 -344 25 -325
rect -25 -361 -17 -344
rect 17 -361 25 -344
rect -25 -369 25 -361
<< polycont >>
rect -17 344 17 361
rect -17 -361 17 -344
<< locali >>
rect -115 413 -67 430
rect 67 413 115 430
rect -115 382 -98 413
rect 98 382 115 413
rect -25 344 -17 361
rect 17 344 25 361
rect -48 319 -31 327
rect -48 -327 -31 -319
rect 31 319 48 327
rect 31 -327 48 -319
rect -25 -361 -17 -344
rect 17 -361 25 -344
rect -115 -413 -98 -382
rect 98 -413 115 -382
rect -115 -430 -67 -413
rect 67 -430 115 -413
<< viali >>
rect -17 344 17 361
rect -48 -319 -31 319
rect 31 -319 48 319
rect -17 -361 17 -344
<< metal1 >>
rect -23 361 23 364
rect -23 344 -17 361
rect 17 344 23 361
rect -23 341 23 344
rect -51 319 -28 325
rect -51 -319 -48 319
rect -31 -319 -28 319
rect -51 -325 -28 -319
rect 28 319 51 325
rect 28 -319 31 319
rect 48 -319 51 319
rect 28 -325 51 -319
rect -23 -344 23 -341
rect -23 -361 -17 -344
rect 17 -361 23 -344
rect -23 -364 23 -361
<< properties >>
string FIXED_BBOX -106 -421 106 421
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 6.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
