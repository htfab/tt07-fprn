magic
tech sky130A
magscale 1 2
timestamp 1717243342
<< locali >>
rect 67 999 246 1195
rect 175 875 342 950
rect 154 426 362 515
rect 77 270 246 376
<< metal1 >>
rect 57 1185 266 1195
rect 57 1100 80 1185
rect 245 1100 266 1185
rect 57 999 266 1100
rect 350 1185 424 1195
rect 350 1100 360 1185
rect 414 1100 424 1185
rect 350 999 424 1100
rect 155 950 362 960
rect 155 875 175 950
rect 342 875 362 950
rect 155 865 362 875
rect 154 505 362 515
rect 154 426 174 505
rect 342 426 362 505
rect 154 416 362 426
rect 57 325 266 386
rect 57 270 77 325
rect 256 270 266 325
rect 57 260 266 270
rect 350 325 424 386
rect 350 270 360 325
rect 414 270 424 325
rect 350 260 424 270
<< via1 >>
rect 80 1100 245 1185
rect 360 1100 414 1185
rect 175 875 342 950
rect 174 426 342 505
rect 77 270 256 325
rect 360 270 414 325
<< metal2 >>
rect 55 1185 255 1290
rect 55 1100 80 1185
rect 245 1100 255 1185
rect 55 1090 255 1100
rect 350 1185 539 1195
rect 350 1100 360 1185
rect 414 1100 539 1185
rect 350 1090 539 1100
rect 154 950 362 960
rect 154 875 175 950
rect 342 875 362 950
rect 154 865 362 875
rect 154 790 255 865
rect 424 790 539 1090
rect 55 590 255 790
rect 340 590 540 790
rect 154 515 255 590
rect 154 505 362 515
rect 154 426 174 505
rect 342 426 362 505
rect 154 416 362 426
rect 424 335 539 590
rect 55 325 266 335
rect 55 270 77 325
rect 256 270 266 325
rect 55 260 266 270
rect 350 325 539 335
rect 350 270 360 325
rect 414 270 539 325
rect 350 260 539 270
rect 55 135 255 260
use sky130_fd_pr__nfet_g5v0d10v5_CYDA8L  XM1
timestamp 1717224314
transform 1 0 308 0 1 323
box -278 -323 278 323
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM2
timestamp 1717224314
transform 1 0 308 0 1 1097
box -308 -397 308 397
<< labels >>
flabel metal2 55 590 255 790 0 FreeSans 256 0 0 0 IN
port 2 nsew
flabel metal2 55 1090 255 1290 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal2 55 135 255 335 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal2 340 590 540 790 0 FreeSans 256 0 0 0 OUT
port 3 nsew
<< end >>
