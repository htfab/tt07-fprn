magic
tech sky130A
magscale 1 2
timestamp 1717244011
<< metal1 >>
rect 1130 13910 30315 14110
rect 4334 13265 4534 13271
rect 4334 13059 4534 13065
rect 9775 11295 9975 13910
rect 14504 13265 14704 13271
rect 14504 13059 14704 13065
rect 19945 11295 20145 13910
rect 24674 13265 24874 13271
rect 24674 13059 24874 13065
rect 30115 11295 30315 13910
rect 9769 11095 9775 11295
rect 9975 11095 9981 11295
rect 19939 11095 19945 11295
rect 20145 11095 20151 11295
rect 30109 11095 30115 11295
rect 30315 11095 30321 11295
<< via1 >>
rect 4334 13065 4534 13265
rect 14504 13065 14704 13265
rect 24674 13065 24874 13265
rect 9775 11095 9975 11295
rect 19945 11095 20145 11295
rect 30115 11095 30315 11295
<< metal2 >>
rect 4339 14110 4529 14114
rect 14509 14110 14699 14114
rect 24679 14110 24869 14114
rect 4335 14105 24873 14110
rect 4335 13915 4339 14105
rect 4529 13915 14509 14105
rect 14699 13915 24679 14105
rect 24869 13915 24873 14105
rect 4335 13910 24873 13915
rect 4339 13906 4529 13910
rect 14509 13906 14699 13910
rect 24679 13906 24869 13910
rect 4334 13435 4534 13444
rect 14504 13435 14704 13444
rect 24674 13435 24874 13444
rect 4328 13065 4334 13265
rect 4534 13065 4540 13265
rect 8912 13024 11210 13245
rect 14498 13065 14504 13265
rect 14704 13065 14710 13265
rect 19082 13024 21380 13245
rect 24668 13065 24674 13265
rect 24874 13065 24880 13265
rect 9775 11295 9975 11301
rect 9775 11089 9975 11095
rect 19945 11295 20145 11301
rect 19945 11089 20145 11095
rect 30115 11295 30315 11301
rect 30115 11089 30315 11095
rect 8910 9864 10386 10087
rect 19080 9864 20556 10087
rect 8912 8509 10385 8730
rect 19082 8509 20555 8730
rect 9756 6580 9765 6780
rect 9965 6580 9974 6780
rect 19926 6580 19935 6780
rect 20135 6580 20144 6780
rect 9115 5349 10411 5572
rect 19285 5349 20581 5572
rect 8779 3810 10391 4031
rect 18949 3810 20561 4031
rect 9110 834 10396 1057
rect 19280 834 20566 1057
<< via2 >>
rect 4339 13915 4529 14105
rect 14509 13915 14699 14105
rect 24679 13915 24869 14105
rect 4334 13265 4534 13435
rect 14504 13265 14704 13435
rect 24674 13265 24874 13435
rect 4334 13235 4534 13265
rect 14504 13235 14704 13265
rect 24674 13235 24874 13265
rect 9765 6580 9965 6780
rect 19935 6580 20135 6780
<< metal3 >>
rect 4334 14105 4534 14110
rect 4334 13915 4339 14105
rect 4529 13915 4534 14105
rect 4334 13440 4534 13915
rect 14504 14105 14704 14110
rect 14504 13915 14509 14105
rect 14699 13915 14704 14105
rect 14504 13440 14704 13915
rect 24674 14105 24874 14110
rect 24674 13915 24679 14105
rect 24869 13915 24874 14105
rect 24674 13440 24874 13915
rect 4329 13435 4539 13440
rect 4329 13235 4334 13435
rect 4534 13235 4539 13435
rect 4329 13230 4539 13235
rect 14499 13435 14709 13440
rect 14499 13235 14504 13435
rect 14704 13235 14709 13435
rect 14499 13230 14709 13235
rect 24669 13435 24879 13440
rect 24669 13235 24674 13435
rect 24874 13235 24879 13435
rect 24669 13230 24879 13235
rect 9760 6780 9970 6785
rect 19930 6780 20140 6785
rect 9760 6580 9765 6780
rect 9965 6580 10380 6780
rect 9760 6575 9970 6580
rect 10180 200 10380 6580
rect 19930 6580 19935 6780
rect 20135 6580 20550 6780
rect 19930 6575 20140 6580
rect 20350 200 20550 6580
rect 10180 0 14635 200
rect 20350 0 24805 200
use grid_cell_ext  grid_cell_ext_0
timestamp 1717244011
transform 1 0 0 0 1 0
box 0 0 9975 13800
use grid_cell_ext  grid_cell_ext_1
timestamp 1717244011
transform 1 0 10170 0 1 0
box 0 0 9975 13800
use grid_cell_ext  grid_cell_ext_2
timestamp 1717244011
transform 1 0 20340 0 1 0
box 0 0 9975 13800
<< end >>
