* NGSPICE file created from inverter.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_CYDA8L a_n108_n65# a_n50_n153# a_n242_n287# a_50_n65#
X0 a_50_n65# a_n50_n153# a_n108_n65# a_n242_n287# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1885 pd=1.88 as=0.1885 ps=1.88 w=0.65 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLAZY6 a_n50_n197# a_50_n100# w_n308_n397# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt inverter VDD IN OUT VSS
XXM1 VSS IN VSS OUT sky130_fd_pr__nfet_g5v0d10v5_CYDA8L
XXM2 IN OUT VDD VDD sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
.ends

