magic
tech sky130A
magscale 1 2
timestamp 1717244011
<< metal2 >>
rect 29740 42910 29930 42914
rect 23935 42905 29935 42910
rect 23935 42715 29740 42905
rect 29930 42715 29935 42905
rect 23935 42710 29935 42715
rect 29740 42706 29930 42710
rect 29331 39900 29340 40090
rect 29530 39900 29539 40090
rect 30935 35580 31135 35589
rect 29960 35380 30935 35580
rect 30935 35371 31135 35380
rect 19570 28505 19760 28514
rect 19570 28306 19760 28315
rect 19161 25500 19170 25690
rect 19360 25500 19369 25690
rect 30535 21180 30735 21189
rect 29985 20980 30535 21180
rect 30535 20971 30735 20980
rect 9400 14105 9590 14114
rect 9400 13906 9590 13915
rect 8991 11100 9000 11290
rect 9190 11100 9199 11290
rect 30135 6780 30335 6789
rect 29995 6580 30135 6780
rect 30135 6571 30335 6580
<< via2 >>
rect 29740 42715 29930 42905
rect 29340 39900 29530 40090
rect 30935 35380 31135 35580
rect 19570 28315 19760 28505
rect 19170 25500 19360 25690
rect 30535 20980 30735 21180
rect 9400 13915 9590 14105
rect 9000 11100 9190 11290
rect 30135 6580 30335 6780
<< metal3 >>
rect 29736 42910 29934 42915
rect 29735 42909 29935 42910
rect 29735 42711 29736 42909
rect 29934 42711 29935 42909
rect 29735 42710 29935 42711
rect 29736 42705 29934 42710
rect 29335 40094 29535 40095
rect 29330 39896 29336 40094
rect 29534 39896 29540 40094
rect 29335 39895 29535 39896
rect 30930 35585 31140 35591
rect 30930 35380 30935 35385
rect 31135 35380 31140 35385
rect 30930 35375 31140 35380
rect 3911 29000 4109 29005
rect 3910 28999 4465 29000
rect 3910 28801 3911 28999
rect 4109 28801 4465 28999
rect 3910 28800 4465 28801
rect 14081 28999 14279 29005
rect 3911 28795 4109 28800
rect 14081 28795 14279 28801
rect 24251 28999 24449 29005
rect 24251 28795 24449 28801
rect 19566 28510 19764 28515
rect 19565 28509 19765 28510
rect 19565 28311 19566 28509
rect 19764 28311 19765 28509
rect 19565 28310 19765 28311
rect 19566 28305 19764 28310
rect 19165 25694 19365 25695
rect 19160 25496 19166 25694
rect 19364 25496 19370 25694
rect 19165 25495 19365 25496
rect 30530 21185 30740 21191
rect 30530 20980 30535 20985
rect 30735 20980 30740 20985
rect 30530 20975 30740 20980
rect 3911 14600 4109 14605
rect 3910 14599 4465 14600
rect 3910 14401 3911 14599
rect 4109 14401 4465 14599
rect 3910 14400 4465 14401
rect 14081 14599 14279 14605
rect 3911 14395 4109 14400
rect 14081 14395 14279 14401
rect 24251 14599 24449 14605
rect 24251 14395 24449 14401
rect 9396 14110 9594 14115
rect 9395 14109 9595 14110
rect 9395 13911 9396 14109
rect 9594 13911 9595 14109
rect 9395 13910 9595 13911
rect 9396 13905 9594 13910
rect 8995 11294 9195 11295
rect 8990 11096 8996 11294
rect 9194 11096 9200 11294
rect 8995 11095 9195 11096
rect 30130 6785 30340 6791
rect 30130 6580 30135 6585
rect 30335 6580 30340 6585
rect 30130 6575 30340 6580
rect 9355 0 9555 200
<< via3 >>
rect 29736 42905 29934 42909
rect 29736 42715 29740 42905
rect 29740 42715 29930 42905
rect 29930 42715 29934 42905
rect 29736 42711 29934 42715
rect 29336 40090 29534 40094
rect 29336 39900 29340 40090
rect 29340 39900 29530 40090
rect 29530 39900 29534 40090
rect 29336 39896 29534 39900
rect 30930 35580 31140 35585
rect 30930 35385 30935 35580
rect 30935 35385 31135 35580
rect 31135 35385 31140 35580
rect 3911 28801 4109 28999
rect 14081 28801 14279 28999
rect 24251 28801 24449 28999
rect 19566 28505 19764 28509
rect 19566 28315 19570 28505
rect 19570 28315 19760 28505
rect 19760 28315 19764 28505
rect 19566 28311 19764 28315
rect 19166 25690 19364 25694
rect 19166 25500 19170 25690
rect 19170 25500 19360 25690
rect 19360 25500 19364 25690
rect 19166 25496 19364 25500
rect 30530 21180 30740 21185
rect 30530 20985 30535 21180
rect 30535 20985 30735 21180
rect 30735 20985 30740 21180
rect 3911 14401 4109 14599
rect 14081 14401 14279 14599
rect 24251 14401 24449 14599
rect 9396 14105 9594 14109
rect 9396 13915 9400 14105
rect 9400 13915 9590 14105
rect 9590 13915 9594 14105
rect 9396 13911 9594 13915
rect 8996 11290 9194 11294
rect 8996 11100 9000 11290
rect 9000 11100 9190 11290
rect 9190 11100 9194 11290
rect 8996 11096 9194 11100
rect 30130 6780 30340 6785
rect 30130 6585 30135 6780
rect 30135 6585 30335 6780
rect 30335 6585 30340 6780
<< metal4 >>
rect 145 307 465 42910
rect 785 307 985 42910
rect 1185 307 1385 42910
rect 1585 307 1785 42910
rect 2285 307 2605 42910
rect 3910 29570 4110 42910
rect 3910 28999 4110 29000
rect 3910 28801 3911 28999
rect 4109 28801 4110 28999
rect 3910 15170 4110 28801
rect 3910 14599 4110 14600
rect 3910 14401 3911 14599
rect 4109 14401 4110 14599
rect 3910 308 4110 14401
rect 4310 308 4510 42910
rect 4710 308 4910 42910
rect 5230 307 5550 42910
rect 5870 307 6070 42910
rect 6270 307 6470 42910
rect 6670 307 6870 42910
rect 7370 307 7690 42910
rect 8995 11294 9195 42910
rect 8995 11096 8996 11294
rect 9194 11096 9195 11294
rect 8995 308 9195 11096
rect 9395 14109 9595 42910
rect 9395 13911 9396 14109
rect 9594 13911 9595 14109
rect 9395 308 9595 13911
rect 10315 307 10635 42910
rect 10955 307 11155 42910
rect 11355 307 11555 42910
rect 11755 307 11955 42910
rect 12455 307 12775 42910
rect 14080 29570 14280 42910
rect 14080 28999 14280 29000
rect 14080 28801 14081 28999
rect 14279 28801 14280 28999
rect 14080 15170 14280 28801
rect 14080 14599 14280 14600
rect 14080 14401 14081 14599
rect 14279 14401 14280 14599
rect 14080 308 14280 14401
rect 14480 308 14680 42910
rect 14880 308 15080 42910
rect 15400 307 15720 42910
rect 16040 307 16240 42910
rect 16440 307 16640 42910
rect 16840 307 17040 42910
rect 17540 307 17860 42910
rect 19165 25694 19365 42910
rect 19165 25496 19166 25694
rect 19364 25496 19365 25694
rect 19165 308 19365 25496
rect 19565 28509 19765 42910
rect 19565 28311 19566 28509
rect 19764 28311 19765 28509
rect 19565 308 19765 28311
rect 20485 307 20805 42910
rect 21125 307 21325 42910
rect 21525 307 21725 42910
rect 21925 307 22125 42910
rect 22625 307 22945 42910
rect 24250 29570 24450 42910
rect 24250 28999 24450 29000
rect 24250 28801 24251 28999
rect 24449 28801 24450 28999
rect 24250 15170 24450 28801
rect 24250 14599 24450 14600
rect 24250 14401 24251 14599
rect 24449 14401 24450 14599
rect 24250 308 24450 14401
rect 24650 308 24850 42910
rect 25050 308 25250 42910
rect 25570 307 25890 42910
rect 26210 307 26410 42910
rect 26610 307 26810 42910
rect 27010 307 27210 42910
rect 27710 307 28030 42910
rect 29335 40094 29535 42910
rect 29335 39896 29336 40094
rect 29534 39896 29535 40094
rect 29335 308 29535 39896
rect 29735 42909 29935 42915
rect 29735 42711 29736 42909
rect 29934 42711 29935 42909
rect 29735 308 29935 42711
rect 30135 6786 30335 42911
rect 30535 21186 30735 42911
rect 30935 35586 31135 42911
rect 30929 35585 31141 35586
rect 30929 35385 30930 35585
rect 31140 35385 31141 35585
rect 30929 35384 31141 35385
rect 30529 21185 30741 21186
rect 30529 20985 30530 21185
rect 30740 20985 30741 21185
rect 30529 20984 30741 20985
rect 30129 6785 30341 6786
rect 30129 6585 30130 6785
rect 30340 6585 30341 6785
rect 30129 6584 30341 6585
rect 30135 308 30335 6584
rect 30535 307 30735 20984
rect 30935 307 31135 35384
use mini_grid_row  mini_grid_row_0
timestamp 1717244011
transform 1 0 0 0 1 0
box 0 0 30321 14114
use mini_grid_row  mini_grid_row_1
timestamp 1717244011
transform 1 0 0 0 1 14400
box 0 0 30321 14114
use mini_grid_row  mini_grid_row_2
timestamp 1717244011
transform 1 0 0 0 1 28800
box 0 0 30321 14114
<< labels >>
flabel metal4 2285 42590 2605 42910 0 FreeSans 240 0 0 0 VSS
port 27 nsew
flabel metal3 9355 0 9555 200 0 FreeSans 128 0 0 0 ANALOG_PIN
port 20 nsew
flabel metal4 785 42710 985 42910 0 FreeSans 128 0 0 0 VD_RES
port 4 nsew
flabel metal4 1185 42710 1385 42910 0 FreeSans 128 0 0 0 VD_SHORT
port 3 nsew
flabel metal4 1585 42710 1785 42910 0 FreeSans 128 0 0 0 VD_LINE
port 2 nsew
flabel metal4 145 42590 465 42910 0 FreeSans 240 0 0 0 VDD
port 1 nsew
flabel metal4 5230 42590 5550 42910 0 FreeSans 240 0 0 0 VDD
port 1 nsew
flabel metal4 10315 42590 10635 42910 0 FreeSans 240 0 0 0 VDD
port 1 nsew
flabel metal4 15400 42590 15720 42910 0 FreeSans 240 0 0 0 VDD
port 1 nsew
flabel metal4 20485 42590 20805 42910 0 FreeSans 240 0 0 0 VDD
port 1 nsew
flabel metal4 25570 42590 25890 42910 0 FreeSans 240 0 0 0 VDD
port 1 nsew
flabel metal4 7370 42590 7690 42910 0 FreeSans 240 0 0 0 VSS
port 27 nsew
flabel metal4 12455 42590 12775 42910 0 FreeSans 240 0 0 0 VSS
port 27 nsew
flabel metal4 17540 42590 17860 42910 0 FreeSans 240 0 0 0 VSS
port 27 nsew
flabel metal4 22625 42590 22945 42910 0 FreeSans 240 0 0 0 VSS
port 27 nsew
flabel metal4 27710 42590 28030 42910 0 FreeSans 240 0 0 0 VSS
port 27 nsew
flabel metal4 5870 42710 6070 42910 0 FreeSans 128 0 0 0 HD_RES
port 7 nsew
flabel metal4 6270 42710 6470 42910 0 FreeSans 128 0 0 0 HD_SHORT
port 6 nsew
flabel metal4 6670 42710 6870 42910 0 FreeSans 128 0 0 0 HD_LINE
port 5 nsew
flabel metal4 16840 42710 17040 42910 0 FreeSans 128 0 0 0 HD_LINE
port 5 nsew
flabel metal4 16440 42710 16640 42910 0 FreeSans 128 0 0 0 HD_SHORT
port 6 nsew
flabel metal4 16040 42710 16240 42910 0 FreeSans 128 0 0 0 HD_RES
port 7 nsew
flabel metal4 11755 42710 11955 42910 0 FreeSans 128 0 0 0 VD_LINE
port 2 nsew
flabel metal4 11355 42710 11555 42910 0 FreeSans 128 0 0 0 VD_SHORT
port 3 nsew
flabel metal4 10955 42710 11155 42910 0 FreeSans 128 0 0 0 VD_RES
port 4 nsew
flabel metal4 27010 42710 27210 42910 0 FreeSans 128 0 0 0 HD_LINE
port 5 nsew
flabel metal4 26610 42710 26810 42910 0 FreeSans 128 0 0 0 HD_SHORT
port 6 nsew
flabel metal4 26210 42710 26410 42910 0 FreeSans 128 0 0 0 HD_RES
port 7 nsew
flabel metal4 21925 42710 22125 42910 0 FreeSans 128 0 0 0 VD_LINE
port 2 nsew
flabel metal4 21525 42710 21725 42910 0 FreeSans 128 0 0 0 VD_SHORT
port 3 nsew
flabel metal4 21125 42710 21325 42910 0 FreeSans 128 0 0 0 VD_RES
port 4 nsew
flabel metal4 3910 42710 4110 42910 0 FreeSans 128 0 0 0 V_INPUT_0
port 14 nsew
flabel metal4 4710 42710 4910 42910 0 FreeSans 128 0 0 0 V_GATE_0
port 8 nsew
flabel metal4 14080 42710 14280 42910 0 FreeSans 128 0 0 0 V_INPUT_1
port 15 nsew
flabel metal4 14880 42710 15080 42910 0 FreeSans 128 0 0 0 V_GATE_1
port 9 nsew
flabel metal4 24250 42710 24450 42910 0 FreeSans 128 0 0 0 V_INPUT_2
port 16 nsew
flabel metal4 25050 42710 25250 42910 0 FreeSans 128 0 0 0 V_GATE_2
port 10 nsew
flabel metal4 4310 42710 4510 42910 0 FreeSans 128 0 0 0 V_LINE_0
port 21 nsew
flabel metal4 14480 42710 14680 42910 0 FreeSans 128 0 0 0 V_LINE_1
port 22 nsew
flabel metal4 24650 42710 24850 42910 0 FreeSans 128 0 0 0 V_LINE_2
port 23 nsew
flabel metal4 8995 42710 9195 42910 0 FreeSans 128 0 0 0 H_LINE_0
port 24 nsew
flabel metal4 9395 42710 9595 42910 0 FreeSans 128 0 0 0 H_GATE_0
port 11 nsew
flabel metal4 19165 42710 19365 42910 0 FreeSans 128 0 0 0 H_LINE_1
port 25 nsew
flabel metal4 19565 42710 19765 42910 0 FreeSans 128 0 0 0 H_GATE_1
port 12 nsew
flabel metal4 29335 42710 29535 42910 0 FreeSans 128 0 0 0 H_LINE_2
port 26 nsew
flabel metal4 29735 42710 29935 42910 0 FreeSans 128 0 0 0 H_GATE_2
port 13 nsew
flabel metal4 30135 42710 30335 42910 0 FreeSans 128 0 0 0 H_INPUT_0
port 17 nsew
flabel metal4 30535 42710 30735 42910 0 FreeSans 128 0 0 0 H_INPUT_1
port 18 nsew
flabel metal4 30935 42710 31135 42910 0 FreeSans 128 0 0 0 H_INPUT_2
port 19 nsew
<< end >>
