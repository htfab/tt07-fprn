magic
tech sky130A
magscale 1 2
timestamp 1717224314
<< pwell >>
rect -201 -1473 201 1473
<< psubdiff >>
rect -165 1403 -69 1437
rect 69 1403 165 1437
rect -165 1341 -131 1403
rect 131 1341 165 1403
rect -165 -1403 -131 -1341
rect 131 -1403 165 -1341
rect -165 -1437 -69 -1403
rect 69 -1437 165 -1403
<< psubdiffcont >>
rect -69 1403 69 1437
rect -165 -1341 -131 1341
rect 131 -1341 165 1341
rect -69 -1437 69 -1403
<< xpolycontact >>
rect -35 875 35 1307
rect -35 -1307 35 -875
<< xpolyres >>
rect -35 -875 35 875
<< locali >>
rect -165 1403 -69 1437
rect 69 1403 165 1437
rect -165 1341 -131 1403
rect 131 1341 165 1403
rect -165 -1403 -131 -1341
rect 131 -1403 165 -1341
rect -165 -1437 -69 -1403
rect 69 -1437 165 -1403
<< viali >>
rect -19 892 19 1289
rect -19 -1289 19 -892
<< metal1 >>
rect -25 1289 25 1301
rect -25 892 -19 1289
rect 19 892 25 1289
rect -25 880 25 892
rect -25 -892 25 -880
rect -25 -1289 -19 -892
rect 19 -1289 25 -892
rect -25 -1301 25 -1289
<< properties >>
string FIXED_BBOX -148 -1420 148 1420
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 8.75 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 51.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
