magic
tech sky130A
magscale 1 2
timestamp 1717243586
<< locali >>
rect 210 4210 410 4300
rect 210 140 410 220
<< viali >>
rect 78 3699 112 3900
rect 504 3699 538 3900
rect 78 539 112 742
rect 504 539 538 742
<< metal1 >>
rect 210 4290 410 4300
rect 210 4220 230 4290
rect 390 4220 410 4290
rect 210 4210 410 4220
rect 58 3900 132 3910
rect 58 3699 68 3900
rect 122 3699 132 3900
rect 58 3689 132 3699
rect 484 3900 558 3910
rect 484 3699 494 3900
rect 548 3699 558 3900
rect 484 3689 558 3699
rect 192 3155 266 3165
rect 192 2179 202 3155
rect 256 2179 266 3155
rect 192 2169 266 2179
rect 350 3155 424 3165
rect 350 2179 360 3155
rect 414 2179 424 3155
rect 350 2169 424 2179
rect 192 1546 266 1556
rect 192 930 202 1546
rect 256 930 266 1546
rect 192 920 266 930
rect 350 1546 424 1556
rect 350 930 360 1546
rect 414 930 424 1546
rect 350 920 424 930
rect 58 742 132 752
rect 58 539 68 742
rect 122 539 132 742
rect 58 529 132 539
rect 484 742 558 752
rect 484 539 494 742
rect 548 539 558 742
rect 484 529 558 539
rect 210 210 410 220
rect 210 150 230 210
rect 390 150 410 210
rect 210 140 410 150
<< via1 >>
rect 230 4220 390 4290
rect 68 3699 78 3900
rect 78 3699 112 3900
rect 112 3699 122 3900
rect 494 3699 504 3900
rect 504 3699 538 3900
rect 538 3699 548 3900
rect 202 2179 256 3155
rect 360 2179 414 3155
rect 202 930 256 1546
rect 360 930 414 1546
rect 68 539 78 742
rect 78 539 112 742
rect 112 539 122 742
rect 494 539 504 742
rect 504 539 538 742
rect 538 539 548 742
rect 230 150 390 210
<< metal2 >>
rect 210 4290 410 4300
rect 210 4220 230 4290
rect 390 4220 410 4290
rect 210 4100 410 4220
rect 58 3900 558 3910
rect 58 3699 68 3900
rect 122 3699 494 3900
rect 548 3699 558 3900
rect 58 3689 558 3699
rect 192 3155 266 3165
rect 192 2179 202 3155
rect 256 2179 266 3155
rect 192 1960 266 2179
rect 65 1760 266 1960
rect 192 1546 266 1760
rect 192 930 202 1546
rect 256 930 266 1546
rect 192 920 266 930
rect 350 3155 424 3165
rect 350 2179 360 3155
rect 414 2179 424 3155
rect 350 1960 424 2179
rect 350 1760 550 1960
rect 350 1546 424 1760
rect 350 930 360 1546
rect 414 930 424 1546
rect 350 920 424 930
rect 58 742 558 752
rect 58 539 68 742
rect 122 539 494 742
rect 548 539 558 742
rect 58 529 558 539
rect 210 210 410 340
rect 210 150 230 210
rect 390 150 410 210
rect 210 140 410 150
use sky130_fd_pr__nfet_g5v0d10v5_TMGAGH  XM1
timestamp 1717243586
transform 1 0 308 0 1 908
box -278 -908 278 908
use sky130_fd_pr__pfet_g5v0d10v5_KLP5N5  XM2
timestamp 1717224314
transform 1 0 308 0 1 3167
box -308 -1297 308 1297
<< labels >>
flabel metal2 210 140 410 340 0 FreeSans 256 0 0 0 EN
port 5 nsew
flabel metal2 210 4100 410 4300 0 FreeSans 256 0 0 0 ENB
port 2 nsew
flabel metal2 65 1760 265 1960 0 FreeSans 256 0 0 0 UA
port 3 nsew
flabel metal2 350 1760 550 1960 0 FreeSans 256 0 0 0 UB
port 4 nsew
flabel metal2 210 540 410 740 0 FreeSans 256 0 0 0 VSS
port 6 nsew
flabel metal2 210 3700 410 3900 0 FreeSans 256 0 0 0 VDD
port 1 nsew
<< end >>
