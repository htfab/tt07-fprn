magic
tech sky130A
magscale 1 2
timestamp 1717244011
<< nwell >>
rect 4112 12700 4135 13494
<< metal1 >>
rect 4340 12755 4540 12955
rect 4885 12755 5085 12955
rect 4600 11925 4821 11931
rect 4600 10997 4821 11704
rect 4600 10776 5722 10997
<< via1 >>
rect 4600 11704 4821 11925
<< metal2 >>
rect 3995 13295 6130 13495
rect 3995 12925 4195 13295
rect 5090 13090 5470 13295
rect 3704 12725 4195 12925
rect 5546 12590 5555 12790
rect 5755 12590 5764 12790
rect 5930 12730 6130 13295
rect 2871 12563 3071 12572
rect 3710 12563 3900 12567
rect 3071 12558 3905 12563
rect 3071 12368 3710 12558
rect 3900 12368 3905 12558
rect 3071 12363 3905 12368
rect 2871 12354 3071 12363
rect 3710 12359 3900 12363
rect 5110 12135 5470 12335
rect 4600 11926 4821 11935
rect 4591 11705 4600 11926
rect 4821 11705 4830 11926
rect 4594 11704 4600 11705
rect 4821 11704 4827 11705
rect 4695 10790 4895 10990
rect 5110 9782 5310 12135
rect 9780 10790 9980 10990
rect 3689 9565 5310 9782
rect 3689 9559 5309 9565
rect 3690 8204 5315 8425
rect 4685 6275 4885 6475
rect 9770 6275 9970 6475
rect 3689 5044 5309 5267
rect 15 3700 215 3900
rect 3700 3726 3921 3910
rect 5091 3726 5312 3910
rect 3700 3505 5312 3726
rect 15 540 215 740
rect 3689 529 5309 752
<< via2 >>
rect 5555 12590 5755 12790
rect 2871 12363 3071 12563
rect 3710 12368 3900 12558
rect 4600 11925 4821 11926
rect 4600 11705 4821 11925
<< metal3 >>
rect 5258 12790 5770 12800
rect 5258 12590 5555 12790
rect 5755 12590 5770 12790
rect 5258 12579 5770 12590
rect 2866 12563 3076 12568
rect 2866 12465 2871 12563
rect 2526 12363 2871 12465
rect 3071 12363 3076 12563
rect 2526 12265 3076 12363
rect 3705 12558 3905 12563
rect 3705 12368 3710 12558
rect 3900 12368 3905 12558
rect 5258 12434 5479 12579
rect 3705 11926 3905 12368
rect 4599 12213 5479 12434
rect 4599 11931 4820 12213
rect 4595 11926 4826 11931
rect 3705 11715 4600 11926
rect 3710 11705 4600 11715
rect 4821 11705 4826 11926
rect 4595 11700 4826 11705
rect 850 9950 1050 10150
rect 5935 9950 6135 10150
rect 850 5435 1050 5635
rect 5935 5435 6135 5635
rect 850 920 1050 1120
rect 4270 -105 4470 1560
rect 5935 920 6135 1120
rect 9361 -105 9561 1560
rect 4270 -305 9561 -105
use resistor_cell  x1
timestamp 1717243805
transform 1 0 -404 0 1 0
box 410 0 5300 13494
use resistor_cell  x2
timestamp 1717243805
transform 1 0 4681 0 1 0
box 410 0 5300 13494
use and_gate  x3
timestamp 1717244011
transform 1 0 4135 0 1 12000
box 0 0 1696 1494
<< labels >>
flabel metal3 4270 -305 4470 -105 0 FreeSans 256 0 0 0 NODE
port 14 nsew
flabel metal3 850 920 1050 1120 0 FreeSans 256 0 0 0 VD_RES
port 8 nsew
flabel metal3 850 5435 1050 5635 0 FreeSans 256 0 0 0 VD_SHORT
port 7 nsew
flabel metal3 850 9950 1050 10150 0 FreeSans 256 0 0 0 VD_LINE
port 5 nsew
flabel metal2 4685 6275 4885 6475 0 FreeSans 256 0 0 0 V_NEXT
port 6 nsew
flabel metal2 4695 10790 4895 10990 0 FreeSans 256 0 0 0 V_LINE
port 4 nsew
flabel metal1 4340 12755 4540 12955 0 FreeSans 256 0 0 0 H_GATE
port 2 nsew
flabel metal1 4885 12755 5085 12955 0 FreeSans 256 0 0 0 V_GATE
port 3 nsew
flabel metal2 15 540 215 740 0 FreeSans 256 0 0 0 VSS
port 15 nsew
flabel metal2 15 3700 215 3900 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal3 5935 920 6135 1120 0 FreeSans 256 0 0 0 HD_RES
port 13 nsew
flabel metal3 5935 5435 6135 5635 0 FreeSans 256 0 0 0 HD_SHORT
port 12 nsew
flabel metal3 5935 9950 6135 10150 0 FreeSans 256 0 0 0 HD_LINE
port 10 nsew
flabel metal2 9780 10790 9980 10990 0 FreeSans 256 0 0 0 H_LINE
port 9 nsew
flabel metal2 9770 6275 9970 6475 0 FreeSans 256 0 0 0 H_NEXT
port 11 nsew
<< end >>
