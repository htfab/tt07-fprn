magic
tech sky130A
magscale 1 2
timestamp 1717249730
<< metal1 >>
rect 7040 45060 7240 45066
rect 17210 45060 17410 45066
rect 27380 45060 27580 45066
rect 512 44860 7040 45060
rect 7240 44860 17210 45060
rect 17410 44860 27380 45060
rect 27580 44860 31509 45060
rect 7040 44854 7240 44860
rect 17210 44854 17410 44860
rect 27380 44854 27580 44860
rect 6640 44710 6840 44716
rect 16810 44710 17010 44716
rect 26980 44710 27180 44716
rect 512 44510 6640 44710
rect 6840 44510 16810 44710
rect 17010 44510 26980 44710
rect 27180 44510 31509 44710
rect 6640 44504 6840 44510
rect 16810 44504 17010 44510
rect 26980 44504 27180 44510
rect 6240 44360 6440 44366
rect 16410 44360 16610 44366
rect 26580 44360 26780 44366
rect 512 44160 6240 44360
rect 6440 44160 16410 44360
rect 16610 44160 26580 44360
rect 26780 44160 31509 44360
rect 6240 44154 6440 44160
rect 16410 44154 16610 44160
rect 26580 44154 26780 44160
rect 1955 44010 2155 44016
rect 12125 44010 12325 44016
rect 22295 44010 22495 44016
rect 25755 44010 25955 44016
rect 512 43810 1955 44010
rect 2155 43810 12125 44010
rect 12325 43810 22295 44010
rect 22495 43810 25755 44010
rect 25955 43810 31509 44010
rect 1955 43804 2155 43810
rect 12125 43804 12325 43810
rect 22295 43804 22495 43810
rect 25755 43804 25955 43810
rect 1555 43660 1755 43666
rect 11725 43660 11925 43666
rect 21895 43660 22095 43666
rect 25015 43660 25215 43666
rect 512 43460 1555 43660
rect 1755 43460 11725 43660
rect 11925 43460 21895 43660
rect 22095 43460 25015 43660
rect 25215 43460 31509 43660
rect 1555 43454 1755 43460
rect 11725 43454 11925 43460
rect 21895 43454 22095 43460
rect 25015 43454 25215 43460
rect 1155 43310 1355 43316
rect 11325 43310 11525 43316
rect 21495 43310 21695 43316
rect 24285 43310 24485 43316
rect 516 43110 1155 43310
rect 1355 43110 11325 43310
rect 11525 43110 21495 43310
rect 21695 43110 24285 43310
rect 24485 43110 31509 43310
rect 1155 43104 1355 43110
rect 11325 43104 11525 43110
rect 21495 43104 21695 43110
rect 24285 43104 24485 43110
<< via1 >>
rect 7040 44860 7240 45060
rect 17210 44860 17410 45060
rect 27380 44860 27580 45060
rect 6640 44510 6840 44710
rect 16810 44510 17010 44710
rect 26980 44510 27180 44710
rect 6240 44160 6440 44360
rect 16410 44160 16610 44360
rect 26580 44160 26780 44360
rect 1955 43810 2155 44010
rect 12125 43810 12325 44010
rect 22295 43810 22495 44010
rect 25755 43810 25955 44010
rect 1555 43460 1755 43660
rect 11725 43460 11925 43660
rect 21895 43460 22095 43660
rect 25015 43460 25215 43660
rect 1155 43110 1355 43310
rect 11325 43110 11525 43310
rect 21495 43110 21695 43310
rect 24285 43110 24485 43310
<< metal2 >>
rect 27960 45060 28160 45069
rect 7034 44860 7040 45060
rect 7240 44860 7246 45060
rect 17204 44860 17210 45060
rect 17410 44860 17416 45060
rect 27374 44860 27380 45060
rect 27580 44860 27960 45060
rect 28160 44860 28169 45060
rect 6634 44510 6640 44710
rect 6840 44510 6846 44710
rect 6234 44160 6240 44360
rect 6440 44160 6446 44360
rect 1949 43810 1955 44010
rect 2155 43810 2161 44010
rect 1546 43460 1555 43660
rect 1755 43460 1764 43660
rect 1160 43310 1350 43314
rect 1149 43110 1155 43310
rect 1355 43110 1361 43310
rect 1555 43304 1755 43460
rect 1555 43114 1560 43304
rect 1750 43114 1755 43304
rect 1160 43106 1350 43110
rect 1555 43109 1755 43114
rect 1955 43305 2155 43810
rect 1955 43115 1960 43305
rect 2150 43115 2155 43305
rect 1955 43110 2155 43115
rect 6240 43305 6440 44160
rect 6240 43115 6245 43305
rect 6435 43115 6440 43305
rect 6240 43110 6440 43115
rect 6640 43305 6840 44510
rect 6640 43115 6645 43305
rect 6835 43115 6840 43305
rect 6640 43110 6840 43115
rect 7040 43305 7240 44860
rect 16804 44510 16810 44710
rect 17010 44510 17016 44710
rect 16404 44160 16410 44360
rect 16610 44160 16616 44360
rect 12119 43810 12125 44010
rect 12325 43810 12331 44010
rect 11716 43460 11725 43660
rect 11925 43460 11934 43660
rect 11330 43310 11520 43314
rect 7040 43115 7045 43305
rect 7235 43115 7240 43305
rect 7040 43110 7240 43115
rect 11319 43110 11325 43310
rect 11525 43110 11531 43310
rect 11725 43304 11925 43460
rect 11725 43114 11730 43304
rect 11920 43114 11925 43304
rect 1560 43105 1750 43109
rect 1960 43106 2150 43110
rect 6245 43106 6435 43110
rect 6645 43106 6835 43110
rect 7045 43106 7235 43110
rect 11330 43106 11520 43110
rect 11725 43109 11925 43114
rect 12125 43305 12325 43810
rect 12125 43115 12130 43305
rect 12320 43115 12325 43305
rect 12125 43110 12325 43115
rect 16410 43305 16610 44160
rect 16410 43115 16415 43305
rect 16605 43115 16610 43305
rect 16410 43110 16610 43115
rect 16810 43305 17010 44510
rect 16810 43115 16815 43305
rect 17005 43115 17010 43305
rect 16810 43110 17010 43115
rect 17210 43305 17410 44860
rect 26980 44710 27180 44719
rect 26974 44510 26980 44710
rect 27180 44510 27186 44710
rect 24285 44360 24485 44369
rect 22289 43810 22295 44010
rect 22495 43810 22501 44010
rect 21886 43460 21895 43660
rect 22095 43460 22104 43660
rect 21500 43310 21690 43314
rect 17210 43115 17215 43305
rect 17405 43115 17410 43305
rect 17210 43110 17410 43115
rect 21489 43110 21495 43310
rect 21695 43110 21701 43310
rect 21895 43304 22095 43460
rect 21895 43114 21900 43304
rect 22090 43114 22095 43304
rect 11730 43105 11920 43109
rect 12130 43106 12320 43110
rect 16415 43106 16605 43110
rect 16815 43106 17005 43110
rect 17215 43106 17405 43110
rect 21500 43106 21690 43110
rect 21895 43109 22095 43114
rect 22295 43305 22495 43810
rect 24285 43310 24485 44160
rect 25015 44360 25215 44369
rect 25015 43660 25215 44160
rect 25755 44360 25955 44369
rect 26580 44360 26780 44369
rect 26574 44160 26580 44360
rect 26780 44160 26786 44360
rect 25755 44010 25955 44160
rect 25749 43810 25755 44010
rect 25955 43810 25961 44010
rect 25009 43460 25015 43660
rect 25215 43460 25221 43660
rect 22295 43115 22300 43305
rect 22490 43115 22495 43305
rect 22295 43110 22495 43115
rect 24279 43110 24285 43310
rect 24485 43110 24491 43310
rect 26580 43305 26780 44160
rect 26580 43115 26585 43305
rect 26775 43115 26780 43305
rect 26580 43110 26780 43115
rect 26980 43305 27180 44510
rect 26980 43115 26985 43305
rect 27175 43115 27180 43305
rect 26980 43110 27180 43115
rect 27380 43305 27580 44860
rect 27960 44851 28160 44860
rect 27380 43115 27385 43305
rect 27575 43115 27580 43305
rect 27380 43110 27580 43115
rect 21900 43105 22090 43109
rect 22300 43106 22490 43110
rect 26585 43106 26775 43110
rect 26985 43106 27175 43110
rect 27385 43106 27575 43110
rect 31287 190 31457 194
rect 9736 185 31462 190
rect 9736 15 31287 185
rect 31457 15 31462 185
rect 9736 10 31462 15
rect 31287 6 31457 10
<< via2 >>
rect 27960 44860 28160 45060
rect 1160 43115 1350 43305
rect 1560 43114 1750 43304
rect 1960 43115 2150 43305
rect 6245 43115 6435 43305
rect 6645 43115 6835 43305
rect 7045 43115 7235 43305
rect 11330 43115 11520 43305
rect 11730 43114 11920 43304
rect 12130 43115 12320 43305
rect 16415 43115 16605 43305
rect 16815 43115 17005 43305
rect 26980 44510 27180 44710
rect 24285 44160 24485 44360
rect 17215 43115 17405 43305
rect 21500 43115 21690 43305
rect 21900 43114 22090 43304
rect 25015 44160 25215 44360
rect 25755 44160 25955 44360
rect 26580 44160 26780 44360
rect 22300 43115 22490 43305
rect 26585 43115 26775 43305
rect 26985 43115 27175 43305
rect 27385 43115 27575 43305
rect 31287 15 31457 185
<< metal3 >>
rect 19130 45060 19330 45066
rect 4280 44860 18395 45060
rect 18595 44860 18601 45060
rect 1156 43310 1354 43315
rect 1155 43309 1355 43310
rect 1556 43309 1754 43314
rect 1956 43310 2154 43315
rect 1955 43309 2155 43310
rect 1155 43111 1156 43309
rect 1354 43111 1355 43309
rect 1155 43110 1355 43111
rect 1555 43308 1755 43309
rect 1555 43110 1556 43308
rect 1754 43110 1755 43308
rect 1955 43111 1956 43309
rect 2154 43111 2155 43309
rect 1955 43110 2155 43111
rect 4280 43309 4480 44860
rect 19130 44710 19330 44860
rect 5080 44510 19330 44710
rect 19860 45060 20060 45066
rect 5080 43309 5280 44510
rect 19860 44360 20060 44860
rect 9765 44160 20060 44360
rect 20600 45060 20800 45066
rect 6641 43310 6839 43315
rect 7041 43310 7239 43315
rect 6240 43309 6440 43310
rect 6640 43309 6840 43310
rect 4280 43111 4281 43309
rect 4479 43111 4480 43309
rect 5075 43111 5081 43309
rect 5279 43111 5285 43309
rect 6235 43111 6241 43309
rect 6439 43111 6445 43309
rect 6640 43111 6641 43309
rect 6839 43111 6840 43309
rect 4280 43110 4480 43111
rect 5080 43110 5280 43111
rect 6240 43110 6440 43111
rect 6640 43110 6840 43111
rect 7040 43309 7240 43310
rect 9765 43309 9965 44160
rect 20600 44010 20800 44860
rect 14450 43810 20800 44010
rect 21335 45060 21535 45066
rect 11326 43310 11524 43315
rect 11325 43309 11525 43310
rect 11726 43309 11924 43314
rect 12126 43310 12324 43315
rect 12125 43309 12325 43310
rect 14450 43309 14650 43810
rect 21335 43660 21535 44860
rect 15250 43460 21535 43660
rect 22075 45060 22275 45066
rect 22075 43659 22275 44860
rect 22075 43461 22076 43659
rect 22274 43461 22275 43659
rect 22075 43460 22275 43461
rect 22810 45060 23010 45066
rect 22810 43660 23010 44860
rect 23545 45060 23745 45066
rect 23545 44010 23745 44860
rect 24285 45060 24485 45066
rect 24285 44365 24485 44860
rect 25015 45060 25215 45066
rect 25015 44365 25215 44860
rect 25755 45060 25955 45066
rect 25755 44365 25955 44860
rect 26490 45060 26690 45066
rect 26490 44365 26690 44860
rect 27225 45060 27425 45066
rect 27225 44715 27425 44860
rect 27955 45065 28165 45071
rect 27955 44849 28165 44855
rect 28695 45060 28895 45066
rect 26975 44710 27425 44715
rect 26975 44510 26980 44710
rect 27180 44510 27425 44710
rect 26975 44505 27185 44510
rect 24280 44360 24490 44365
rect 24280 44160 24285 44360
rect 24485 44160 24490 44360
rect 24280 44155 24490 44160
rect 25010 44360 25220 44365
rect 25010 44160 25015 44360
rect 25215 44160 25220 44360
rect 25010 44155 25220 44160
rect 25750 44360 25960 44365
rect 25750 44160 25755 44360
rect 25955 44160 25960 44360
rect 26490 44360 26785 44365
rect 26490 44160 26580 44360
rect 26780 44160 26785 44360
rect 25750 44155 25960 44160
rect 26575 44155 26785 44160
rect 23545 43810 25620 44010
rect 22810 43460 24820 43660
rect 15250 43309 15450 43460
rect 22076 43455 22274 43460
rect 16811 43310 17009 43315
rect 17211 43310 17409 43315
rect 21496 43310 21694 43315
rect 16410 43309 16610 43310
rect 16810 43309 17010 43310
rect 7040 43111 7041 43309
rect 7239 43111 7240 43309
rect 9760 43111 9766 43309
rect 9964 43111 9970 43309
rect 11325 43111 11326 43309
rect 11524 43111 11525 43309
rect 7040 43110 7240 43111
rect 9765 43110 9965 43111
rect 11325 43110 11525 43111
rect 11725 43308 11925 43309
rect 11725 43110 11726 43308
rect 11924 43110 11925 43308
rect 12125 43111 12126 43309
rect 12324 43111 12325 43309
rect 14445 43111 14451 43309
rect 14649 43111 14655 43309
rect 15245 43111 15251 43309
rect 15449 43111 15455 43309
rect 16405 43111 16411 43309
rect 16609 43111 16615 43309
rect 16810 43111 16811 43309
rect 17009 43111 17010 43309
rect 12125 43110 12325 43111
rect 14450 43110 14650 43111
rect 15250 43110 15450 43111
rect 16410 43110 16610 43111
rect 16810 43110 17010 43111
rect 17210 43309 17410 43310
rect 17210 43111 17211 43309
rect 17409 43111 17410 43309
rect 17210 43110 17410 43111
rect 21495 43309 21695 43310
rect 21896 43309 22094 43314
rect 22296 43310 22494 43315
rect 24620 43314 24820 43460
rect 22295 43309 22495 43310
rect 21495 43111 21496 43309
rect 21694 43111 21695 43309
rect 21495 43110 21695 43111
rect 21895 43308 22095 43309
rect 21895 43110 21896 43308
rect 22094 43110 22095 43308
rect 22295 43111 22296 43309
rect 22494 43111 22495 43309
rect 24615 43116 24621 43314
rect 24819 43116 24825 43314
rect 25420 43309 25620 43810
rect 26981 43310 27179 43315
rect 27381 43310 27579 43315
rect 28695 43310 28895 44860
rect 29430 45060 29630 45066
rect 29430 43660 29630 44860
rect 30170 45060 30370 45066
rect 30170 44010 30370 44860
rect 30900 45060 31100 45066
rect 30900 44360 31100 44860
rect 30900 44160 31505 44360
rect 30170 43810 31105 44010
rect 29430 43460 30705 43660
rect 26580 43309 26780 43310
rect 26980 43309 27180 43310
rect 24620 43115 24820 43116
rect 25415 43111 25421 43309
rect 25619 43111 25625 43309
rect 26575 43111 26581 43309
rect 26779 43111 26785 43309
rect 26980 43111 26981 43309
rect 27179 43111 27180 43309
rect 22295 43110 22495 43111
rect 25420 43110 25620 43111
rect 26580 43110 26780 43111
rect 26980 43110 27180 43111
rect 27380 43309 27580 43310
rect 27380 43111 27381 43309
rect 27579 43111 27580 43309
rect 27380 43110 27580 43111
rect 28695 43309 30305 43310
rect 30505 43309 30705 43460
rect 30905 43309 31105 43810
rect 31305 43309 31505 44160
rect 28695 43111 30106 43309
rect 30304 43111 30310 43309
rect 30500 43111 30506 43309
rect 30704 43111 30710 43309
rect 30900 43111 30906 43309
rect 31104 43111 31110 43309
rect 31300 43111 31306 43309
rect 31504 43111 31510 43309
rect 28695 43110 30305 43111
rect 30505 43110 30705 43111
rect 30905 43110 31105 43111
rect 31305 43110 31505 43111
rect 1156 43105 1354 43110
rect 1555 43109 1755 43110
rect 1556 43104 1754 43109
rect 1956 43105 2154 43110
rect 4281 43105 4479 43110
rect 6641 43105 6839 43110
rect 7041 43105 7239 43110
rect 11326 43105 11524 43110
rect 11725 43109 11925 43110
rect 11726 43104 11924 43109
rect 12126 43105 12324 43110
rect 16811 43105 17009 43110
rect 17211 43105 17409 43110
rect 21496 43105 21694 43110
rect 21895 43109 22095 43110
rect 21896 43104 22094 43109
rect 22296 43105 22494 43110
rect 26981 43105 27179 43110
rect 27381 43105 27579 43110
rect 9715 0 9915 200
rect 31283 190 31461 195
rect 31282 189 31462 190
rect 31282 11 31283 189
rect 31461 11 31462 189
rect 31282 10 31462 11
rect 31283 5 31461 10
<< via3 >>
rect 18395 44860 18595 45060
rect 19130 44860 19330 45060
rect 1156 43305 1354 43309
rect 1156 43115 1160 43305
rect 1160 43115 1350 43305
rect 1350 43115 1354 43305
rect 1156 43111 1354 43115
rect 1556 43304 1754 43308
rect 1556 43114 1560 43304
rect 1560 43114 1750 43304
rect 1750 43114 1754 43304
rect 1556 43110 1754 43114
rect 1956 43305 2154 43309
rect 1956 43115 1960 43305
rect 1960 43115 2150 43305
rect 2150 43115 2154 43305
rect 1956 43111 2154 43115
rect 19860 44860 20060 45060
rect 20600 44860 20800 45060
rect 4281 43111 4479 43309
rect 5081 43111 5279 43309
rect 6241 43305 6439 43309
rect 6241 43115 6245 43305
rect 6245 43115 6435 43305
rect 6435 43115 6439 43305
rect 6241 43111 6439 43115
rect 6641 43305 6839 43309
rect 6641 43115 6645 43305
rect 6645 43115 6835 43305
rect 6835 43115 6839 43305
rect 6641 43111 6839 43115
rect 21335 44860 21535 45060
rect 22075 44860 22275 45060
rect 22076 43461 22274 43659
rect 22810 44860 23010 45060
rect 23545 44860 23745 45060
rect 24285 44860 24485 45060
rect 25015 44860 25215 45060
rect 25755 44860 25955 45060
rect 26490 44860 26690 45060
rect 27225 44860 27425 45060
rect 27955 45060 28165 45065
rect 27955 44860 27960 45060
rect 27960 44860 28160 45060
rect 28160 44860 28165 45060
rect 27955 44855 28165 44860
rect 28695 44860 28895 45060
rect 7041 43305 7239 43309
rect 7041 43115 7045 43305
rect 7045 43115 7235 43305
rect 7235 43115 7239 43305
rect 7041 43111 7239 43115
rect 9766 43111 9964 43309
rect 11326 43305 11524 43309
rect 11326 43115 11330 43305
rect 11330 43115 11520 43305
rect 11520 43115 11524 43305
rect 11326 43111 11524 43115
rect 11726 43304 11924 43308
rect 11726 43114 11730 43304
rect 11730 43114 11920 43304
rect 11920 43114 11924 43304
rect 11726 43110 11924 43114
rect 12126 43305 12324 43309
rect 12126 43115 12130 43305
rect 12130 43115 12320 43305
rect 12320 43115 12324 43305
rect 12126 43111 12324 43115
rect 14451 43111 14649 43309
rect 15251 43111 15449 43309
rect 16411 43305 16609 43309
rect 16411 43115 16415 43305
rect 16415 43115 16605 43305
rect 16605 43115 16609 43305
rect 16411 43111 16609 43115
rect 16811 43305 17009 43309
rect 16811 43115 16815 43305
rect 16815 43115 17005 43305
rect 17005 43115 17009 43305
rect 16811 43111 17009 43115
rect 17211 43305 17409 43309
rect 17211 43115 17215 43305
rect 17215 43115 17405 43305
rect 17405 43115 17409 43305
rect 17211 43111 17409 43115
rect 21496 43305 21694 43309
rect 21496 43115 21500 43305
rect 21500 43115 21690 43305
rect 21690 43115 21694 43305
rect 21496 43111 21694 43115
rect 21896 43304 22094 43308
rect 21896 43114 21900 43304
rect 21900 43114 22090 43304
rect 22090 43114 22094 43304
rect 21896 43110 22094 43114
rect 22296 43305 22494 43309
rect 22296 43115 22300 43305
rect 22300 43115 22490 43305
rect 22490 43115 22494 43305
rect 22296 43111 22494 43115
rect 24621 43116 24819 43314
rect 29430 44860 29630 45060
rect 30170 44860 30370 45060
rect 30900 44860 31100 45060
rect 25421 43111 25619 43309
rect 26581 43305 26779 43309
rect 26581 43115 26585 43305
rect 26585 43115 26775 43305
rect 26775 43115 26779 43305
rect 26581 43111 26779 43115
rect 26981 43305 27179 43309
rect 26981 43115 26985 43305
rect 26985 43115 27175 43305
rect 27175 43115 27179 43305
rect 26981 43111 27179 43115
rect 27381 43305 27579 43309
rect 27381 43115 27385 43305
rect 27385 43115 27575 43305
rect 27575 43115 27579 43305
rect 27381 43111 27579 43115
rect 30106 43111 30304 43309
rect 30506 43111 30704 43309
rect 30906 43111 31104 43309
rect 31306 43111 31504 43309
rect 31283 185 31461 189
rect 31283 15 31287 185
rect 31287 15 31457 185
rect 31457 15 31461 185
rect 31283 11 31461 15
<< metal4 >>
rect 798 44715 858 45152
rect 1534 44715 1594 45152
rect 2270 44715 2330 45152
rect 3006 44715 3066 45152
rect 3742 44715 3802 45152
rect 4478 44715 4538 45152
rect 5214 44715 5274 45152
rect 5950 44715 6010 45152
rect 6686 44715 6746 45152
rect 7422 44715 7482 45152
rect 8158 44715 8218 45152
rect 8894 44715 8954 45152
rect 9630 44715 9690 45152
rect 10366 44715 10426 45152
rect 11102 44715 11162 45152
rect 11838 44715 11898 45152
rect 12574 44715 12634 45152
rect 13310 44715 13370 45152
rect 14046 44715 14106 45152
rect 14782 44715 14842 45152
rect 15518 44715 15578 45152
rect 16254 44715 16314 45152
rect 16990 44715 17050 45152
rect 17726 44715 17786 45152
rect 18462 45061 18522 45152
rect 19198 45061 19258 45152
rect 19934 45061 19994 45152
rect 20670 45061 20730 45152
rect 21406 45061 21466 45152
rect 22142 45061 22202 45152
rect 22878 45061 22938 45152
rect 23614 45061 23674 45152
rect 24350 45061 24410 45152
rect 25086 45061 25146 45152
rect 25822 45061 25882 45152
rect 26558 45061 26618 45152
rect 27294 45061 27354 45152
rect 28030 45066 28090 45152
rect 27954 45065 28166 45066
rect 18394 45060 18596 45061
rect 18394 44860 18395 45060
rect 18595 44860 18596 45060
rect 18394 44859 18596 44860
rect 19129 45060 19331 45061
rect 19129 44860 19130 45060
rect 19330 44860 19331 45060
rect 19129 44859 19331 44860
rect 19859 45060 20061 45061
rect 19859 44860 19860 45060
rect 20060 44860 20061 45060
rect 19859 44859 20061 44860
rect 20599 45060 20801 45061
rect 20599 44860 20600 45060
rect 20800 44860 20801 45060
rect 20599 44859 20801 44860
rect 21334 45060 21536 45061
rect 21334 44860 21335 45060
rect 21535 44860 21536 45060
rect 21334 44859 21536 44860
rect 22074 45060 22276 45061
rect 22074 44860 22075 45060
rect 22275 44860 22276 45060
rect 22074 44859 22276 44860
rect 22809 45060 23011 45061
rect 22809 44860 22810 45060
rect 23010 44860 23011 45060
rect 22809 44859 23011 44860
rect 23544 45060 23746 45061
rect 23544 44860 23545 45060
rect 23745 44860 23746 45060
rect 23544 44859 23746 44860
rect 24284 45060 24486 45061
rect 24284 44860 24285 45060
rect 24485 44860 24486 45060
rect 24284 44859 24486 44860
rect 25014 45060 25216 45061
rect 25014 44860 25015 45060
rect 25215 44860 25216 45060
rect 25014 44859 25216 44860
rect 25754 45060 25956 45061
rect 25754 44860 25755 45060
rect 25955 44860 25956 45060
rect 25754 44859 25956 44860
rect 26489 45060 26691 45061
rect 26489 44860 26490 45060
rect 26690 44860 26691 45060
rect 26489 44859 26691 44860
rect 27224 45060 27426 45061
rect 27224 44860 27225 45060
rect 27425 44860 27426 45060
rect 27224 44859 27426 44860
rect 27954 44855 27955 45065
rect 28165 44855 28166 45065
rect 28766 45061 28826 45152
rect 29502 45061 29562 45152
rect 30238 45061 30298 45152
rect 30974 45061 31034 45152
rect 28694 45060 28896 45061
rect 28694 44860 28695 45060
rect 28895 44860 28896 45060
rect 28694 44859 28896 44860
rect 29429 45060 29631 45061
rect 29429 44860 29430 45060
rect 29630 44860 29631 45060
rect 29429 44859 29631 44860
rect 30169 45060 30371 45061
rect 30169 44860 30170 45060
rect 30370 44860 30371 45060
rect 30169 44859 30371 44860
rect 30899 45060 31101 45061
rect 30899 44860 30900 45060
rect 31100 44860 31101 45060
rect 31710 44952 31770 45152
rect 30899 44859 31101 44860
rect 27954 44854 28166 44855
rect 510 44395 17920 44715
rect 515 307 835 43310
rect 1155 43309 1355 43310
rect 1955 43309 2155 43310
rect 1155 43111 1156 43309
rect 1354 43111 1355 43309
rect 1155 42910 1355 43111
rect 1555 43308 1755 43309
rect 1555 43110 1556 43308
rect 1754 43110 1755 43308
rect 1555 42910 1755 43110
rect 1955 43111 1956 43309
rect 2154 43111 2155 43309
rect 1955 42910 2155 43111
rect 2655 307 2975 44395
rect 19935 43659 22275 43660
rect 19935 43461 22076 43659
rect 22274 43461 22275 43659
rect 19935 43460 22275 43461
rect 4280 43309 4480 43310
rect 4280 43111 4281 43309
rect 4479 43111 4480 43309
rect 4280 42710 4480 43111
rect 5080 43309 5280 43310
rect 5080 43111 5081 43309
rect 5279 43111 5280 43309
rect 5080 42710 5280 43111
rect 5600 307 5920 43310
rect 6240 43309 6440 43310
rect 6240 43111 6241 43309
rect 6439 43111 6440 43309
rect 6240 42910 6440 43111
rect 6640 43309 6840 43310
rect 6640 43111 6641 43309
rect 6839 43111 6840 43309
rect 6640 42910 6840 43111
rect 7040 43309 7240 43310
rect 7040 43111 7041 43309
rect 7239 43111 7240 43309
rect 7040 42910 7240 43111
rect 7740 307 8060 43310
rect 9765 43309 9965 43310
rect 9765 43111 9766 43309
rect 9964 43111 9965 43309
rect 9765 42710 9965 43111
rect 10685 307 11005 43310
rect 11325 43309 11525 43310
rect 12125 43309 12325 43310
rect 11325 43111 11326 43309
rect 11524 43111 11525 43309
rect 11325 42910 11525 43111
rect 11725 43308 11925 43309
rect 11725 43110 11726 43308
rect 11924 43110 11925 43308
rect 11725 42910 11925 43110
rect 12125 43111 12126 43309
rect 12324 43111 12325 43309
rect 12125 42910 12325 43111
rect 12825 307 13145 43310
rect 14450 43309 14650 43310
rect 14450 43111 14451 43309
rect 14649 43111 14650 43309
rect 14450 42710 14650 43111
rect 15250 43309 15450 43310
rect 15250 43111 15251 43309
rect 15449 43111 15450 43309
rect 15250 42710 15450 43111
rect 15770 307 16090 43310
rect 16410 43309 16610 43310
rect 16410 43111 16411 43309
rect 16609 43111 16610 43309
rect 16410 42910 16610 43111
rect 16810 43309 17010 43310
rect 16810 43111 16811 43309
rect 17009 43111 17010 43309
rect 16810 42910 17010 43111
rect 17210 43309 17410 43310
rect 17210 43111 17211 43309
rect 17409 43111 17410 43309
rect 17210 42910 17410 43111
rect 17910 307 18230 43310
rect 19935 42710 20135 43460
rect 24620 43314 24820 43315
rect 20855 307 21175 43310
rect 21495 43309 21695 43310
rect 22295 43309 22495 43310
rect 21495 43111 21496 43309
rect 21694 43111 21695 43309
rect 21495 42910 21695 43111
rect 21895 43308 22095 43309
rect 21895 43110 21896 43308
rect 22094 43110 22095 43308
rect 21895 42910 22095 43110
rect 22295 43111 22296 43309
rect 22494 43111 22495 43309
rect 22295 42910 22495 43111
rect 22995 307 23315 43310
rect 24620 43116 24621 43314
rect 24819 43116 24820 43314
rect 24620 42710 24820 43116
rect 25420 43309 25620 43310
rect 25420 43111 25421 43309
rect 25619 43111 25620 43309
rect 25420 42710 25620 43111
rect 25940 307 26260 43310
rect 26580 43309 26780 43310
rect 26580 43111 26581 43309
rect 26779 43111 26780 43309
rect 26580 42910 26780 43111
rect 26980 43309 27180 43310
rect 26980 43111 26981 43309
rect 27179 43111 27180 43309
rect 26980 42910 27180 43111
rect 27380 43309 27580 43310
rect 27380 43111 27381 43309
rect 27579 43111 27580 43309
rect 27380 42910 27580 43111
rect 28080 307 28400 43310
rect 30105 43309 30305 43310
rect 30105 43111 30106 43309
rect 30304 43111 30305 43309
rect 30105 42710 30305 43111
rect 30505 43309 30705 43310
rect 30505 43111 30506 43309
rect 30704 43111 30705 43309
rect 30505 42711 30705 43111
rect 30905 43309 31105 43310
rect 30905 43111 30906 43309
rect 31104 43111 31105 43309
rect 30905 42711 31105 43111
rect 31305 43309 31505 43310
rect 31305 43111 31306 43309
rect 31504 43111 31505 43309
rect 31305 42711 31505 43111
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 189 31462 200
rect 31282 11 31283 189
rect 31461 11 31462 189
rect 31282 0 31462 11
use mini_grid  mini_grid_0
timestamp 1717244011
transform 1 0 370 0 1 0
box 0 0 31141 42915
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 28080 307 28400 43310 1 FreeSans 800 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 22995 307 23315 43310 1 FreeSans 800 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 17910 307 18230 43310 1 FreeSans 800 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 12825 307 13145 43310 1 FreeSans 800 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 7740 307 8060 43310 1 FreeSans 800 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 2655 307 2975 43310 1 FreeSans 800 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 25940 307 26260 43310 1 FreeSans 800 90 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 20855 307 21175 43310 1 FreeSans 800 90 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 15770 307 16090 43310 1 FreeSans 800 90 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 10685 307 11005 43310 1 FreeSans 800 90 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 5600 307 5920 43310 1 FreeSans 800 90 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 515 307 835 43310 1 FreeSans 800 90 0 0 VPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
