magic
tech sky130A
magscale 1 2
timestamp 1717243586
<< metal1 >>
rect 645 4300 845 4306
rect 1380 4300 1580 4306
rect 845 4100 1030 4300
rect 645 4094 1030 4100
rect 505 3890 705 3900
rect 505 3715 560 3890
rect 695 3715 705 3890
rect 505 2750 705 3715
rect 830 3080 1030 4094
rect 1190 4100 1380 4300
rect 1190 4094 1580 4100
rect 1190 3435 1390 4094
rect 1190 3229 1390 3235
rect 1535 3890 1735 3900
rect 1535 3715 1545 3890
rect 1675 3715 1735 3890
rect 830 2880 1190 3080
rect 1390 2880 1396 3080
rect 1535 2750 1735 3715
rect 505 2740 1735 2750
rect 505 2560 605 2740
rect 785 2560 1145 2740
rect 1325 2560 1735 2740
rect 505 2550 1735 2560
<< via1 >>
rect 645 4100 845 4300
rect 560 3715 695 3890
rect 1380 4100 1580 4300
rect 1190 3235 1390 3435
rect 1545 3715 1675 3890
rect 1190 2880 1390 3080
rect 605 2560 785 2740
rect 1145 2560 1325 2740
<< metal2 >>
rect 210 4100 645 4300
rect 845 4100 851 4300
rect 55 3890 705 3910
rect 1015 3905 1215 4300
rect 1374 4100 1380 4300
rect 1580 4100 2030 4300
rect 55 3715 560 3890
rect 695 3715 705 3890
rect 55 3690 705 3715
rect 830 3705 1215 3905
rect 1535 3890 2180 3910
rect 1535 3715 1545 3890
rect 1675 3715 2180 3890
rect 830 3430 1030 3705
rect 1535 3690 2180 3715
rect 1750 3689 2180 3690
rect 826 3240 835 3430
rect 1025 3240 1034 3430
rect 830 3235 1030 3240
rect 1181 3235 1190 3435
rect 1390 3235 1399 3435
rect 1190 3080 1390 3086
rect 1390 2880 1535 3080
rect 1735 2880 1744 3080
rect 1190 2874 1390 2880
rect 595 2740 795 2750
rect 595 2560 605 2740
rect 785 2560 795 2740
rect 595 2260 795 2560
rect 1135 2740 1335 2750
rect 1135 2560 1145 2740
rect 1325 2560 1335 2740
rect 1135 2260 1335 2560
rect 350 1960 550 1969
rect 65 1760 265 1960
rect 550 1955 795 1960
rect 550 1766 799 1955
rect 550 1760 795 1766
rect 871 1760 880 1960
rect 1080 1760 1335 1960
rect 1420 1760 1886 1960
rect 1961 1760 1970 1960
rect 2170 1760 2179 1960
rect 350 1751 550 1760
rect 595 1255 795 1505
rect 1135 1255 1335 1505
rect 595 1055 1335 1255
rect 1450 1120 1650 1129
rect 1686 1120 1886 1760
rect 595 752 795 1055
rect 1650 920 1886 1120
rect 1450 911 1650 920
rect 59 750 1080 752
rect 1370 750 2176 752
rect 59 529 2176 750
rect 210 335 410 340
rect 1450 335 1650 340
rect 1830 335 2030 340
rect 206 145 215 335
rect 405 145 414 335
rect 1446 145 1455 335
rect 1645 145 1654 335
rect 1826 145 1835 335
rect 2025 145 2034 335
rect 210 140 410 145
rect 1450 140 1650 145
rect 1830 140 2030 145
<< via2 >>
rect 835 3240 1025 3430
rect 1190 3235 1390 3435
rect 1535 2880 1735 3080
rect 350 1760 550 1960
rect 880 1760 1080 1960
rect 1970 1760 2170 1960
rect 1450 920 1650 1120
rect 215 145 405 335
rect 1455 145 1645 335
rect 1835 145 2025 335
<< metal3 >>
rect 350 3904 1215 3905
rect 350 3705 2169 3904
rect 350 1965 550 3705
rect 1185 3435 1395 3440
rect 765 3430 1030 3435
rect 765 3240 835 3430
rect 1025 3240 1030 3430
rect 765 3235 1030 3240
rect 1185 3235 1190 3435
rect 1390 3235 1395 3435
rect 765 1965 965 3235
rect 1185 3230 1395 3235
rect 345 1960 555 1965
rect 345 1760 350 1960
rect 550 1760 555 1960
rect 765 1960 1085 1965
rect 765 1760 880 1960
rect 1080 1760 1085 1960
rect 345 1755 555 1760
rect 875 1755 1085 1760
rect 1190 1505 1390 3230
rect 1530 3080 1740 3085
rect 1530 2880 1535 3080
rect 1735 2880 1740 3080
rect 1530 2875 1740 2880
rect 210 1305 1390 1505
rect 1535 1505 1735 2875
rect 1970 2824 2169 3705
rect 1970 2676 2170 2824
rect 1971 1965 2170 2676
rect 1965 1960 2175 1965
rect 1965 1760 1970 1960
rect 2170 1760 2175 1960
rect 1965 1755 2175 1760
rect 1535 1305 2030 1505
rect 210 335 410 1305
rect 1445 1120 1655 1125
rect 1445 920 1450 1120
rect 1650 920 1655 1120
rect 1445 915 1655 920
rect 210 145 215 335
rect 405 145 410 335
rect 210 140 410 145
rect 1450 335 1650 915
rect 1450 145 1455 335
rect 1645 145 1650 335
rect 1450 140 1650 145
rect 1830 335 2030 1305
rect 1830 145 1835 335
rect 2025 145 2030 335
rect 1830 140 2030 145
use pass_gate  x1
timestamp 1717243586
transform 1 0 0 0 1 0
box 0 0 616 4464
use pass_gate  x2
timestamp 1717243586
transform 1 0 1620 0 1 0
box 0 0 616 4464
use inverter  x3
timestamp 1717243342
transform 1 0 540 0 1 1170
box 0 0 616 1494
use inverter  x4
timestamp 1717243342
transform 1 0 1080 0 1 1170
box 0 0 616 1494
<< labels >>
flabel metal2 210 540 410 740 0 FreeSans 256 0 0 0 VSS
port 7 nsew
flabel metal2 210 3700 410 3900 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel metal2 210 140 410 340 0 FreeSans 256 0 0 0 GATE
port 6 nsew
flabel metal2 210 4100 410 4300 0 FreeSans 256 0 0 0 GATEB
port 4 nsew
flabel metal2 65 1760 265 1960 0 FreeSans 256 0 0 0 D
port 5 nsew
flabel metal2 1450 140 1650 340 0 FreeSans 256 0 0 0 Q
port 1 nsew
flabel metal2 1015 4100 1215 4300 0 FreeSans 256 0 0 0 QB
port 3 nsew
flabel metal2 1830 540 2030 740 0 FreeSans 256 0 0 0 VSS
port 7 nsew
flabel metal2 1830 3700 2030 3900 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel metal2 1830 4100 2030 4300 0 FreeSans 256 0 0 0 GATE
port 6 nsew
flabel metal2 1830 140 2030 340 0 FreeSans 256 0 0 0 GATEB
port 4 nsew
<< end >>
