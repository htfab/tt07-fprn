* NGSPICE file created from pass_gate.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_TMGAGH a_n50_n738# a_50_n650# a_n242_n872# a_n108_n650#
X0 a_50_n650# a_n50_n738# a_n108_n650# a_n242_n872# sky130_fd_pr__nfet_g5v0d10v5 ad=1.885 pd=13.58 as=1.885 ps=13.58 w=6.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLP5N5 a_n108_n1000# a_n50_n1097# a_50_n1000#
+ w_n308_n1297#
X0 a_50_n1000# a_n50_n1097# a_n108_n1000# w_n308_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
.ends

.subckt pass_gate VDD ENB UA UB EN VSS
XXM1 EN UB VSS UA sky130_fd_pr__nfet_g5v0d10v5_TMGAGH
XXM2 UA ENB UB VDD sky130_fd_pr__pfet_g5v0d10v5_KLP5N5
.ends

