magic
tech sky130A
magscale 1 2
timestamp 1717243586
<< metal2 >>
rect 755 4295 945 4304
rect 755 4096 945 4105
rect 1546 4100 1555 4300
rect 1755 4100 1764 4300
rect 2915 4295 3105 4304
rect 2915 4096 3105 4105
rect 50 3690 1100 3910
rect 2215 3690 3260 3910
rect 50 3689 930 3690
rect 50 2260 250 3689
rect 340 1960 540 1969
rect 51 1765 60 1955
rect 250 1765 259 1955
rect 340 1751 540 1760
rect 55 752 255 1505
rect 606 1120 806 1960
rect 2765 1760 2965 1960
rect 3050 1760 3250 1960
rect 366 920 375 1120
rect 575 920 806 1120
rect 54 750 930 752
rect 54 530 1100 750
rect 2210 530 3255 750
rect 54 529 930 530
rect 2714 340 3105 344
rect 2713 335 3110 340
rect 2713 145 2714 335
rect 2904 145 3110 335
rect 2713 140 3110 145
rect 2714 136 3105 140
<< via2 >>
rect 755 4105 945 4295
rect 1555 4100 1755 4300
rect 2915 4105 3105 4295
rect 60 1765 250 1955
rect 340 1760 540 1960
rect 375 920 575 1120
rect 755 145 945 335
rect 1995 145 2185 335
rect 2714 145 2904 335
<< metal3 >>
rect 1550 4300 1760 4305
rect 340 4295 950 4300
rect 340 4105 755 4295
rect 945 4105 950 4295
rect 340 4100 950 4105
rect 1550 4100 1555 4300
rect 1755 4295 3110 4300
rect 1755 4105 2915 4295
rect 3105 4105 3110 4295
rect 1755 4100 3110 4105
rect 340 1965 540 4100
rect 1550 4095 1760 4100
rect 335 1960 545 1965
rect 55 1955 255 1960
rect 55 1765 60 1955
rect 250 1765 255 1955
rect 55 1505 255 1765
rect 335 1760 340 1960
rect 540 1760 545 1960
rect 335 1755 545 1760
rect 55 1305 950 1505
rect 370 1120 580 1125
rect 55 920 375 1120
rect 575 920 580 1120
rect 370 915 580 920
rect 750 335 950 1305
rect 2710 340 2908 345
rect 750 145 755 335
rect 945 145 950 335
rect 750 140 950 145
rect 1984 140 1990 340
rect 2190 140 2196 340
rect 2709 339 2909 340
rect 2709 141 2710 339
rect 2908 141 2909 339
rect 2709 140 2909 141
rect 2710 135 2908 140
<< via3 >>
rect 1990 335 2190 340
rect 1990 145 1995 335
rect 1995 145 2185 335
rect 2185 145 2190 335
rect 1990 140 2190 145
rect 2710 335 2908 339
rect 2710 145 2714 335
rect 2714 145 2904 335
rect 2904 145 2908 335
rect 2710 141 2908 145
<< metal4 >>
rect 1989 340 2191 341
rect 1989 140 1990 340
rect 2190 339 2909 340
rect 2190 141 2710 339
rect 2908 141 2909 339
rect 2190 140 2909 141
rect 1989 139 2191 140
use pass_gate  x1
timestamp 1717243586
transform 1 0 2700 0 1 0
box 0 0 616 4464
use latch  x2
timestamp 1717243586
transform 1 0 540 0 1 0
box 0 0 2236 4464
use inverter  x3
timestamp 1717243342
transform 1 0 0 0 1 1170
box 0 0 616 1494
<< labels >>
flabel metal2 50 3700 250 3900 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal2 55 540 255 740 0 FreeSans 256 0 0 0 VSS
port 7 nsew
flabel metal3 55 1760 255 1960 0 FreeSans 256 0 0 0 GATE
port 4 nsew
flabel metal3 55 920 255 1120 0 FreeSans 256 0 0 0 D
port 3 nsew
flabel metal2 2765 1760 2965 1960 0 FreeSans 256 0 0 0 UA
port 6 nsew
flabel metal2 3050 1760 3250 1960 0 FreeSans 256 0 0 0 UB
port 5 nsew
flabel metal4 1990 140 2190 340 0 FreeSans 256 0 0 0 Q
port 2 nsew
<< end >>
