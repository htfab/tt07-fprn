magic
tech sky130A
magscale 1 2
timestamp 1717244011
<< locali >>
rect 90 1010 246 1185
rect 360 994 455 1200
rect 697 994 796 1200
rect 895 1009 1079 1195
rect 210 865 405 955
rect 750 865 945 955
rect 210 430 405 515
rect 274 426 342 430
rect 192 376 266 391
rect 192 270 202 376
rect 256 270 266 376
rect 192 255 266 270
rect 350 376 424 391
rect 350 270 360 376
rect 414 270 424 376
rect 350 255 424 270
rect 504 144 648 502
rect 750 430 945 515
rect 814 426 882 430
rect 732 376 806 391
rect 732 270 742 376
rect 796 270 806 376
rect 732 255 806 270
rect 895 270 910 376
rect 944 366 1079 376
rect 1064 270 1079 366
rect 895 260 1079 270
<< viali >>
rect 202 270 256 376
rect 360 270 414 376
rect 742 270 796 376
rect 910 366 944 376
rect 910 270 1064 366
<< metal1 >>
rect 955 1200 1155 1320
rect 360 1185 796 1200
rect 360 1010 490 1185
rect 660 1010 796 1185
rect 360 994 796 1010
rect 895 1120 1155 1200
rect 895 1009 1079 1120
rect 205 420 405 960
rect 750 420 950 960
rect 142 381 271 391
rect 142 265 152 381
rect 261 265 271 381
rect 142 255 271 265
rect 350 376 806 391
rect 350 270 360 376
rect 414 270 742 376
rect 796 270 806 376
rect 350 255 806 270
rect 895 270 910 376
rect 944 366 1079 376
rect 1064 345 1079 366
rect 1064 270 1155 345
rect 895 260 1155 270
rect 905 255 1155 260
rect 955 145 1155 255
<< via1 >>
rect 490 1010 660 1185
rect 152 376 261 381
rect 152 270 202 376
rect 202 270 256 376
rect 256 270 261 376
rect 152 265 261 270
<< metal2 >>
rect 475 1185 675 1200
rect 475 1010 490 1185
rect 660 1010 675 1185
rect 475 425 675 1010
rect 105 381 675 425
rect 105 265 152 381
rect 261 265 675 381
rect 105 225 675 265
use sky130_fd_pr__nfet_g5v0d10v5_CYDA8L  XM1
timestamp 1717224314
transform 1 0 308 0 1 323
box -278 -323 278 323
use sky130_fd_pr__nfet_g5v0d10v5_CYDA8L  XM2
timestamp 1717224314
transform 1 0 848 0 1 323
box -278 -323 278 323
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM3
timestamp 1717224314
transform 1 0 308 0 1 1097
box -308 -397 308 397
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM4
timestamp 1717224314
transform 1 0 848 0 1 1097
box -308 -397 308 397
<< labels >>
flabel metal1 205 590 405 790 0 FreeSans 256 0 0 0 A
port 2 nsew
flabel metal1 750 590 950 790 0 FreeSans 256 0 0 0 B
port 4 nsew
flabel metal2 475 225 675 425 0 FreeSans 256 0 0 0 OUT
port 3 nsew
flabel metal1 955 145 1155 345 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 955 1120 1155 1320 0 FreeSans 256 0 0 0 VDD
port 1 nsew
<< end >>
