magic
tech sky130A
magscale 1 2
timestamp 1717243805
<< locali >>
rect 4687 4495 4855 4505
rect 4687 4461 4702 4495
rect 4840 4461 4855 4495
rect 4687 4451 4855 4461
rect 4726 3918 4816 4380
rect 4726 2183 4816 2198
rect 4726 1751 4736 2183
rect 4806 1751 4816 2183
rect 4726 1736 4816 1751
rect 4692 1655 4850 1665
rect 4692 1621 4702 1655
rect 4840 1621 4850 1655
rect 4692 1611 4850 1621
<< viali >>
rect 4702 4461 4840 4495
rect 4736 1751 4806 2183
rect 4702 1621 4840 1655
<< metal1 >>
rect 830 10990 1030 11001
rect 824 10790 830 10990
rect 1030 10790 1036 10990
rect 830 10145 1030 10790
rect 420 9945 1030 10145
rect 420 6475 620 9945
rect 821 9781 1044 9792
rect 815 9558 821 9781
rect 1044 9558 1050 9781
rect 414 6275 420 6475
rect 620 6275 626 6475
rect 420 1960 620 6275
rect 821 5266 1044 9558
rect 815 5043 821 5266
rect 1044 5043 1050 5266
rect 4657 5044 4663 5267
rect 4886 5044 4892 5267
rect 414 1760 420 1960
rect 620 1760 626 1960
rect 420 1754 620 1760
rect 821 752 1044 5043
rect 4663 4495 4886 5044
rect 4663 4461 4702 4495
rect 4840 4461 4886 4495
rect 4663 4449 4886 4461
rect 4726 4260 4816 4380
rect 4726 3933 4736 4260
rect 4806 3933 4816 4260
rect 4726 3918 4816 3933
rect 4726 2183 4816 2198
rect 4726 1751 4736 2183
rect 4806 1751 4816 2183
rect 4726 1736 4816 1751
rect 4658 1655 4881 1666
rect 4658 1621 4702 1655
rect 4840 1621 4881 1655
rect 4658 752 4881 1621
rect 812 529 821 752
rect 1044 529 1052 752
rect 821 523 1044 529
rect 4658 523 4881 529
<< via1 >>
rect 830 10790 1030 10990
rect 821 9558 1044 9781
rect 420 6275 620 6475
rect 821 5043 1044 5266
rect 4663 5044 4886 5267
rect 420 1760 620 1960
rect 4736 3933 4806 4260
rect 4736 1751 4806 2183
rect 821 529 1044 752
rect 4658 529 4881 752
<< metal2 >>
rect 1239 12940 1460 12949
rect 1233 12719 1239 12940
rect 1460 12719 1471 12940
rect 1239 12710 1460 12719
rect 830 10995 1030 10996
rect 824 10990 1036 10995
rect 815 10790 830 10990
rect 1030 10985 1455 10990
rect 1030 10795 1260 10985
rect 1450 10795 1455 10985
rect 1030 10790 1455 10795
rect 830 10784 1030 10790
rect 3965 10490 4165 10990
rect 4250 10790 5300 10990
rect 3961 10300 3970 10490
rect 4160 10300 4169 10490
rect 3965 10295 4165 10300
rect 821 9786 1044 9787
rect 815 9782 1050 9786
rect 410 9781 1477 9782
rect 410 9559 821 9781
rect 1044 9559 1477 9781
rect 1044 9558 1336 9559
rect 821 9552 1044 9558
rect 825 8426 1036 8430
rect 755 8425 1240 8426
rect 410 8421 1471 8425
rect 410 8210 825 8421
rect 1036 8210 1471 8421
rect 410 8204 1471 8210
rect 825 8201 1036 8204
rect 420 6480 620 6481
rect 414 6475 626 6480
rect 410 6275 420 6475
rect 620 6470 1455 6475
rect 620 6280 1260 6470
rect 1450 6280 1455 6470
rect 620 6275 1455 6280
rect 420 6269 620 6275
rect 3965 6075 4165 6475
rect 4250 6275 5290 6475
rect 3961 5885 3970 6075
rect 4160 5885 4169 6075
rect 3965 5880 4165 5885
rect 4671 5650 4871 6275
rect 4667 5460 4676 5650
rect 4866 5460 4875 5650
rect 4671 5455 4871 5460
rect 821 5267 1044 5272
rect 4663 5267 4886 5273
rect 410 5266 1477 5267
rect 410 5044 821 5266
rect 815 5043 821 5044
rect 1044 5044 1477 5266
rect 4235 5044 4663 5267
rect 1044 5043 1461 5044
rect 821 5037 1044 5043
rect 4663 5038 4886 5044
rect 4671 4250 4736 4260
rect 4806 4250 4871 4260
rect 4671 4041 4736 4050
rect 4726 3933 4736 4041
rect 4806 4041 4871 4050
rect 4806 3933 4816 4041
rect 4726 3918 4816 3933
rect 620 3910 1460 3911
rect 410 3906 1471 3910
rect 410 3695 825 3906
rect 1036 3695 1471 3906
rect 410 3689 1471 3695
rect 4726 2183 4816 2198
rect 4726 2070 4736 2183
rect 420 1960 620 1966
rect 4670 1960 4736 2070
rect 410 1760 420 1960
rect 620 1955 1455 1960
rect 620 1765 1260 1955
rect 1450 1765 1455 1955
rect 620 1760 1455 1765
rect 420 1754 620 1760
rect 3966 1560 4166 1960
rect 4250 1760 4736 1960
rect 4726 1751 4736 1760
rect 4806 2070 4816 2183
rect 4806 1760 4870 2070
rect 4806 1751 4816 1760
rect 4726 1736 4816 1751
rect 3957 1360 3966 1560
rect 4166 1360 4175 1560
rect 818 752 1046 758
rect 410 529 821 752
rect 1044 529 1477 752
rect 4104 529 4658 752
rect 4881 529 4887 752
rect 818 523 1046 529
<< via2 >>
rect 1239 12719 1460 12940
rect 1260 10795 1450 10985
rect 3970 10300 4160 10490
rect 825 8210 1036 8421
rect 1260 6280 1450 6470
rect 3970 5885 4160 6075
rect 4676 5460 4866 5650
rect 4671 4050 4736 4250
rect 4736 4050 4806 4250
rect 4806 4050 4871 4250
rect 825 3695 1036 3906
rect 1260 1765 1450 1955
rect 3966 1360 4166 1560
<< metal3 >>
rect 1234 12940 1465 12945
rect 1234 12719 1239 12940
rect 1460 12719 1465 12940
rect 1234 12714 1465 12719
rect 1239 12046 1460 12714
rect 820 11825 1460 12046
rect 820 8431 1041 11825
rect 3965 10490 4870 10495
rect 3965 10300 3970 10490
rect 4160 10300 4870 10490
rect 3965 10295 4870 10300
rect 1255 9950 1455 10150
rect 815 8421 1046 8431
rect 815 8210 825 8421
rect 1036 8210 1046 8421
rect 815 8200 1046 8210
rect 820 3916 1041 8200
rect 4670 6080 4870 10295
rect 3965 6075 5290 6080
rect 3965 5885 3970 6075
rect 4160 5885 5290 6075
rect 3965 5880 5290 5885
rect 4671 5650 4871 5655
rect 1255 5435 1455 5635
rect 4671 5460 4676 5650
rect 4866 5460 4871 5650
rect 4671 4255 4871 5460
rect 4666 4250 4876 4255
rect 4666 4050 4671 4250
rect 4871 4050 4876 4250
rect 4666 4045 4876 4050
rect 815 3906 1046 3916
rect 815 3695 825 3906
rect 1036 3695 1046 3906
rect 5090 3810 5290 5880
rect 815 3685 1046 3695
rect 4680 3610 5290 3810
rect 3961 1560 4171 1565
rect 4680 1560 4880 3610
rect 3961 1360 3966 1560
rect 4166 1360 4880 1560
rect 3961 1355 4171 1360
rect 1255 920 1455 1120
use latched_switch  x1
timestamp 1717243586
transform 1 0 1200 0 1 0
box 0 0 3316 4464
use latched_switch  x2
timestamp 1717243586
transform 1 0 1200 0 1 4515
box 0 0 3316 4464
use latched_switch  x3
timestamp 1717243586
transform 1 0 1200 0 1 9030
box 0 0 3316 4464
use sky130_fd_pr__res_xhigh_po_0p35_75WWSS  XR1
timestamp 1717224314
transform 1 0 4771 0 1 3058
box -201 -1473 201 1473
<< labels >>
flabel metal3 1255 920 1455 1120 0 FreeSans 256 0 0 0 D_RES
port 6 nsew
flabel metal3 1255 5435 1455 5635 0 FreeSans 256 0 0 0 D_SHORT
port 4 nsew
flabel metal3 1255 9950 1455 10150 0 FreeSans 256 0 0 0 D_LINE
port 3 nsew
flabel metal3 5090 5880 5290 6080 0 FreeSans 256 0 0 0 UA
port 8 nsew
flabel metal2 5090 6275 5290 6475 0 FreeSans 256 0 0 0 UB
port 5 nsew
flabel metal2 5100 10790 5300 10990 0 FreeSans 256 0 0 0 LINE
port 2 nsew
flabel metal2 420 3700 620 3900 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal2 420 1760 620 1960 0 FreeSans 256 0 0 0 GATE
port 7 nsew
flabel metal2 420 540 620 740 0 FreeSans 256 0 0 0 VSS
port 9 nsew
<< end >>
