magic
tech sky130A
magscale 1 2
timestamp 1717244011
<< metal1 >>
rect 955 1290 1155 1320
rect 925 1090 935 1290
rect 1130 1090 1155 1290
rect 205 590 405 955
rect 750 590 950 955
rect 955 335 1155 345
rect 924 135 930 335
rect 1130 145 1155 335
rect 1130 135 1136 145
<< via1 >>
rect 935 1090 1130 1290
rect 930 135 1130 335
<< metal2 >>
rect 930 1290 1130 1296
rect 930 1090 935 1290
rect 1130 1090 1335 1290
rect 930 1084 1130 1090
rect 1135 610 1335 790
rect 475 410 1335 610
rect 1420 590 1620 790
rect 475 225 675 410
rect 930 335 1130 341
rect 1130 135 1335 335
rect 930 129 1130 135
use nand_gate  x1
timestamp 1717244011
transform 1 0 0 0 1 0
box 0 0 1156 1494
use inverter  x2
timestamp 1717243342
transform 1 0 1080 0 1 0
box 0 0 616 1494
<< labels >>
flabel metal2 1135 1090 1335 1290 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal2 1135 135 1335 335 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 205 755 405 955 0 FreeSans 256 0 0 0 A
port 3 nsew
flabel metal1 750 755 950 955 0 FreeSans 256 0 0 0 B
port 4 nsew
flabel metal2 1420 590 1620 790 0 FreeSans 256 0 0 0 OUT
port 2 nsew
<< end >>
