magic
tech sky130A
magscale 1 2
timestamp 1717244011
<< metal1 >>
rect 4879 13259 5079 13265
rect 4879 13053 5079 13059
<< via1 >>
rect 4879 13059 5079 13259
<< metal2 >>
rect 4879 13259 5079 13268
rect 4873 13059 4879 13259
rect 5079 13059 5085 13259
rect 4879 13050 5079 13059
rect 4315 11291 4505 11300
rect 4315 11092 4505 11101
rect 2345 10075 2545 10087
rect 2345 9866 2545 9875
rect 7430 10075 7630 10087
rect 7430 9866 7630 9875
rect 3840 6776 4105 6785
rect 3840 6586 3915 6776
rect 3840 6577 4105 6586
rect 2345 5560 2545 5572
rect 2345 5351 2545 5360
rect 7430 5560 7630 5572
rect 7430 5351 7630 5360
rect 406 4000 415 4211
rect 626 4000 635 4211
rect 2345 1045 2545 1057
rect 2345 836 2545 845
rect 7430 1045 7630 1057
rect 7430 836 7630 845
<< via2 >>
rect 4879 13059 5079 13259
rect 4315 11101 4505 11291
rect 2345 9875 2545 10075
rect 7430 9875 7630 10075
rect 3915 6586 4105 6776
rect 2345 5360 2545 5560
rect 7430 5360 7630 5560
rect 415 4000 626 4211
rect 2345 845 2545 1045
rect 7430 845 7630 1045
<< metal3 >>
rect 4874 13259 5084 13264
rect 4710 13258 4879 13259
rect 191 13245 414 13251
rect 414 13024 1041 13245
rect 4705 13060 4711 13258
rect 4710 13059 4879 13060
rect 5079 13059 5084 13259
rect 4874 13054 5084 13059
rect 191 13018 414 13024
rect 5276 12351 5499 12357
rect 5499 12130 5715 12351
rect 5276 12124 5499 12130
rect 4311 11296 4509 11301
rect 4310 11295 4510 11296
rect 4310 11097 4311 11295
rect 4509 11097 4510 11295
rect 4310 11096 4510 11097
rect 4311 11091 4509 11096
rect 1165 9400 1365 10454
rect 2340 10080 2550 10086
rect 2340 9875 2345 9880
rect 2545 9875 2550 9880
rect 2340 9870 2550 9875
rect 6250 9400 6450 10454
rect 7425 10080 7635 10086
rect 7425 9875 7430 9880
rect 7630 9875 7635 9880
rect 7425 9870 7635 9875
rect 1165 9399 1785 9400
rect 6250 9399 6870 9400
rect 1165 9201 1586 9399
rect 1784 9201 1790 9399
rect 6250 9201 6671 9399
rect 6869 9201 6875 9399
rect 1165 9200 1785 9201
rect 6250 9200 6870 9201
rect 191 8730 414 8736
rect 191 8503 414 8509
rect 5276 8730 5499 8736
rect 5276 8503 5499 8509
rect 3911 6781 4109 6786
rect 3910 6780 4110 6781
rect 3910 6582 3911 6780
rect 4109 6582 4110 6780
rect 3910 6581 4110 6582
rect 3911 6576 4109 6581
rect 1185 5940 1385 5946
rect 6270 5940 6470 5946
rect 965 5740 1185 5940
rect 6050 5740 6270 5940
rect 1185 5734 1385 5740
rect 6270 5734 6470 5740
rect 2340 5565 2550 5571
rect 2340 5360 2345 5365
rect 2545 5360 2550 5365
rect 2340 5355 2550 5360
rect 7425 5565 7635 5571
rect 7425 5360 7430 5365
rect 7630 5360 7635 5365
rect 7425 5355 7635 5360
rect 410 4216 414 4221
rect 404 3995 410 4216
rect 621 4211 631 4216
rect 626 4000 631 4211
rect 621 3995 631 4000
rect 5276 4215 5499 4221
rect 410 3990 414 3995
rect 5276 3988 5499 3994
rect 846 1425 1044 1430
rect 5931 1425 6129 1430
rect 845 1424 1221 1425
rect 845 1226 846 1424
rect 1044 1226 1221 1424
rect 845 1225 1221 1226
rect 5930 1424 6306 1425
rect 5930 1226 5931 1424
rect 6129 1226 6306 1424
rect 5930 1225 6306 1226
rect 846 1220 1044 1225
rect 5931 1220 6129 1225
rect 2340 1050 2550 1056
rect 2340 845 2345 850
rect 2545 845 2550 850
rect 2340 840 2550 845
rect 7425 1050 7635 1056
rect 7425 845 7430 850
rect 7630 845 7635 850
rect 7425 840 7635 845
<< via3 >>
rect 191 13024 414 13245
rect 4711 13060 4879 13258
rect 4879 13060 4909 13258
rect 5276 12130 5499 12351
rect 4311 11291 4509 11295
rect 4311 11101 4315 11291
rect 4315 11101 4505 11291
rect 4505 11101 4509 11291
rect 4311 11097 4509 11101
rect 2340 10075 2550 10080
rect 2340 9880 2345 10075
rect 2345 9880 2545 10075
rect 2545 9880 2550 10075
rect 7425 10075 7635 10080
rect 7425 9880 7430 10075
rect 7430 9880 7630 10075
rect 7630 9880 7635 10075
rect 1586 9201 1784 9399
rect 6671 9201 6869 9399
rect 191 8509 414 8730
rect 5276 8509 5499 8730
rect 3911 6776 4109 6780
rect 3911 6586 3915 6776
rect 3915 6586 4105 6776
rect 4105 6586 4109 6776
rect 3911 6582 4109 6586
rect 1185 5740 1385 5940
rect 6270 5740 6470 5940
rect 2340 5560 2550 5565
rect 2340 5365 2345 5560
rect 2345 5365 2545 5560
rect 2545 5365 2550 5560
rect 7425 5560 7635 5565
rect 7425 5365 7430 5560
rect 7430 5365 7630 5560
rect 7630 5365 7635 5560
rect 410 4211 621 4216
rect 410 4000 415 4211
rect 415 4000 621 4211
rect 410 3995 621 4000
rect 5276 3994 5499 4215
rect 846 1226 1044 1424
rect 5931 1226 6129 1424
rect 2340 1045 2550 1050
rect 2340 850 2345 1045
rect 2345 850 2545 1045
rect 2545 850 2550 1045
rect 7425 1045 7635 1050
rect 7425 850 7430 1045
rect 7430 850 7630 1045
rect 7630 850 7635 1045
<< metal4 >>
rect 145 13245 465 13352
rect 145 13024 191 13245
rect 414 13024 465 13245
rect 145 8730 465 13024
rect 145 8509 191 8730
rect 414 8509 465 8730
rect 145 4217 465 8509
rect 145 4216 622 4217
rect 145 3995 410 4216
rect 621 3995 622 4216
rect 145 3994 622 3995
rect 145 768 465 3994
rect 785 1425 985 13352
rect 1185 5941 1385 13352
rect 1585 9399 1785 13352
rect 1585 9201 1586 9399
rect 1784 9201 1785 9399
rect 1184 5940 1386 5941
rect 1184 5740 1185 5940
rect 1385 5740 1386 5940
rect 1184 5739 1386 5740
rect 785 1424 1051 1425
rect 785 1226 846 1424
rect 1044 1226 1051 1424
rect 785 1225 1051 1226
rect 785 768 985 1225
rect 1185 768 1385 5739
rect 1585 768 1785 9201
rect 2285 10080 2605 13351
rect 2285 9880 2340 10080
rect 2550 9880 2605 10080
rect 2285 5565 2605 9880
rect 2285 5365 2340 5565
rect 2550 5365 2605 5565
rect 2285 1050 2605 5365
rect 2285 850 2340 1050
rect 2550 850 2605 1050
rect 2285 768 2605 850
rect 3910 6780 4110 13351
rect 3910 6582 3911 6780
rect 4109 6582 4110 6780
rect 3910 770 4110 6582
rect 4310 11295 4510 13351
rect 4310 11097 4311 11295
rect 4509 11097 4510 11295
rect 4310 770 4510 11097
rect 4710 13258 4910 13351
rect 4710 13060 4711 13258
rect 4909 13060 4910 13258
rect 4710 770 4910 13060
rect 5230 12351 5550 13351
rect 5230 12130 5276 12351
rect 5499 12130 5550 12351
rect 5230 8730 5550 12130
rect 5230 8509 5276 8730
rect 5499 8509 5550 8730
rect 5230 4215 5550 8509
rect 5230 3994 5276 4215
rect 5499 3994 5550 4215
rect 5230 770 5550 3994
rect 5870 1425 6070 13351
rect 6270 5941 6470 13351
rect 6670 9399 6870 13351
rect 6670 9201 6671 9399
rect 6869 9201 6870 9399
rect 6269 5940 6471 5941
rect 6269 5740 6270 5940
rect 6470 5740 6471 5940
rect 6269 5739 6471 5740
rect 5870 1424 6136 1425
rect 5870 1226 5931 1424
rect 6129 1226 6136 1424
rect 5870 1225 6136 1226
rect 5870 770 6070 1225
rect 6270 770 6470 5739
rect 6670 770 6870 9201
rect 7370 10080 7690 13351
rect 7370 9880 7425 10080
rect 7635 9880 7690 10080
rect 7370 5565 7690 9880
rect 7370 5365 7425 5565
rect 7635 5365 7690 5565
rect 7370 1050 7690 5365
rect 7370 850 7425 1050
rect 7635 850 7690 1050
rect 7370 768 7690 850
rect 8995 770 9195 13351
rect 9395 770 9595 13351
use grid_cell  x1
timestamp 1717244011
transform 1 0 -6 0 1 305
box 6 -305 9981 13495
<< end >>
